
module huffman_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module huffman_DW01_add_1 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2XL U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module huffman_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
endmodule


module huffman_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_2 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_3 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_4 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_5 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2XL U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVXL U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module huffman_DW01_inc_6 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2XL U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVXL U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module huffman ( clk, reset, gray_valid, gray_data, CNT_valid, CNT1, CNT2, 
        CNT3, CNT4, CNT5, CNT6, code_valid, HC1, HC2, HC3, HC4, HC5, HC6, M1, 
        M2, M3, M4, M5, M6 );
  input [7:0] gray_data;
  output [7:0] CNT1;
  output [7:0] CNT2;
  output [7:0] CNT3;
  output [7:0] CNT4;
  output [7:0] CNT5;
  output [7:0] CNT6;
  output [7:0] HC1;
  output [7:0] HC2;
  output [7:0] HC3;
  output [7:0] HC4;
  output [7:0] HC5;
  output [7:0] HC6;
  output [7:0] M1;
  output [7:0] M2;
  output [7:0] M3;
  output [7:0] M4;
  output [7:0] M5;
  output [7:0] M6;
  input clk, reset, gray_valid;
  output CNT_valid, code_valid;
  wire   n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, \int_k[2] ,
         N296, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387,
         N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398,
         N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409,
         N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420,
         N421, N422, N423, N424, N425, N440, N441, N442, N443, N444, N445,
         N446, \ListA[0][3] , \ListA[0][2] , \ListA[0][1] , \ListA[0][0] ,
         \ListA[1][3] , \ListA[1][2] , \ListA[1][1] , \ListA[1][0] ,
         \ListA[2][3] , \ListA[2][2] , \ListA[2][1] , \ListA[2][0] ,
         \ListA[3][3] , \ListA[3][2] , \ListA[3][1] , \ListA[3][0] ,
         \ListA[4][3] , \ListA[4][2] , \ListA[4][1] , \ListA[4][0] ,
         \ListA[5][3] , \ListA[5][2] , \ListA[5][1] , \ListA[5][0] ,
         \ListB[0][7] , \ListB[0][6] , \ListB[0][5] , \ListB[0][4] ,
         \ListB[0][3] , \ListB[0][2] , \ListB[0][1] , \ListB[0][0] ,
         \ListB[1][7] , \ListB[1][6] , \ListB[1][5] , \ListB[1][4] ,
         \ListB[1][3] , \ListB[1][2] , \ListB[1][1] , \ListB[1][0] ,
         \ListB[2][7] , \ListB[2][6] , \ListB[2][5] , \ListB[2][4] ,
         \ListB[2][3] , \ListB[2][2] , \ListB[2][1] , \ListB[2][0] ,
         \ListB[3][7] , \ListB[3][6] , \ListB[3][5] , \ListB[3][4] ,
         \ListB[3][3] , \ListB[3][2] , \ListB[3][1] , \ListB[3][0] ,
         \ListB[4][7] , \ListB[4][6] , \ListB[4][5] , \ListB[4][4] ,
         \ListB[4][3] , \ListB[4][2] , \ListB[4][1] , \ListB[4][0] ,
         \ListB[5][7] , \ListB[5][6] , \ListB[5][5] , \ListB[5][4] ,
         \ListB[5][3] , \ListB[5][2] , \ListB[5][1] , \ListB[5][0] , N488,
         N492, N493, N494, N495, N496, N497, N498, N499, \Tree_1[1][3] ,
         \Tree_1[1][2] , \Tree_1[1][1] , \Tree_1[1][0] , \Tree_1[2][3] ,
         \Tree_1[2][2] , \Tree_1[2][1] , \Tree_1[2][0] , \Tree_1[4][3] ,
         \Tree_1[4][2] , \Tree_1[4][1] , \Tree_1[4][0] , \Tree_0[1][3] ,
         \Tree_0[1][2] , \Tree_0[1][1] , \Tree_0[1][0] , \Tree_0[2][3] ,
         \Tree_0[2][2] , \Tree_0[2][1] , \Tree_0[2][0] , \Tree_0[4][3] ,
         \Tree_0[4][2] , \Tree_0[4][1] , \Tree_0[4][0] , N712, N713, N714,
         N715, N716, N717, N718, N719, N774, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n139, n140, n149, n150, n151, n246, n247,
         n248, n249, n251, n252, n253, n255, n256, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n309, n310, n311, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n351, n352, n353, n354, n355, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n390, n391, n392, n393, n394, n396, n397, n398, n399,
         n400, n401, n403, n406, n409, n413, n415, n418, n420, n421, n422,
         n424, n425, n426, n428, n429, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n455, n456, n457, n458, n459, n460, n461,
         n462, n470, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n595, n602, n604, n605,
         n606, n608, n609, n611, n612, n613, n615, n616, n618, n619, n620,
         n622, n623, n624, n625, n626, n627, n629, n630, n631, n632, n633,
         n634, n636, n637, n639, n640, n641, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n661, n662, n669, n676, n683, n690, n697, n704, n705, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, net5452, net5500, net5501, net5512, net5660, net5661,
         net5701, net7156, net7189, net7188, net5477, net5475, net7390,
         net7492, net7476, net7469, net7595, n914, n915, n916, n917, n918,
         n919, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, net7494, net7433, net7388, net7385,
         net7366, net5697, net5514, net5488, n933, n932, n931, n1215, n1217,
         n1219, n1221, n1223, n1225, n1227, n1229, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243;
  wire   [2:0] cs;
  wire   [6:0] cnt;
  wire   [2:0] int_j;
  wire   [2:0] int_i;
  wire   [3:0] cnt2;
  wire   [3:0] RegA_t;
  wire   [7:0] RegA_v;
  wire   [7:0] RegB_v;
  wire   [3:0] RegB_t;
  wire   [3:0] node;
  wire   [3:0] tmp_T1;
  wire   [3:0] tmp_T0;
  wire   [7:0] addnum;
  wire   [7:0] tmp_HC;

  DFFRX2 \CNT6_reg[7]  ( .D(n873), .CK(clk), .RN(n1045), .Q(CNT6[7]), .QN(n107) );
  DFFRX2 \CNT6_reg[6]  ( .D(n874), .CK(clk), .RN(n1084), .Q(CNT6[6]), .QN(n108) );
  DFFRX2 \CNT6_reg[5]  ( .D(n875), .CK(clk), .RN(n1045), .Q(CNT6[5]), .QN(n109) );
  DFFRX2 \CNT6_reg[4]  ( .D(n876), .CK(clk), .RN(n1045), .Q(CNT6[4]), .QN(n110) );
  DFFRX2 \CNT6_reg[3]  ( .D(n877), .CK(clk), .RN(n1045), .Q(CNT6[3]), .QN(n111) );
  DFFRX2 \CNT6_reg[2]  ( .D(n878), .CK(clk), .RN(n1045), .Q(CNT6[2]), .QN(n112) );
  DFFRX2 \CNT6_reg[1]  ( .D(n879), .CK(clk), .RN(n1047), .Q(CNT6[1]), .QN(n113) );
  DFFRX2 \CNT6_reg[0]  ( .D(n880), .CK(clk), .RN(n1047), .Q(CNT6[0]), .QN(n114) );
  DFFRX2 \CNT3_reg[7]  ( .D(n881), .CK(clk), .RN(n1047), .Q(CNT3[7]), .QN(n99)
         );
  DFFRX2 \CNT3_reg[6]  ( .D(n882), .CK(clk), .RN(n1047), .Q(CNT3[6]), .QN(n100) );
  DFFRX2 \CNT3_reg[5]  ( .D(n883), .CK(clk), .RN(n1047), .Q(CNT3[5]), .QN(n101) );
  DFFRX2 \CNT3_reg[4]  ( .D(n884), .CK(clk), .RN(n1047), .Q(CNT3[4]), .QN(n102) );
  DFFRX2 \CNT3_reg[3]  ( .D(n885), .CK(clk), .RN(n1047), .Q(CNT3[3]), .QN(n103) );
  DFFRX2 \CNT3_reg[2]  ( .D(n886), .CK(clk), .RN(n1047), .Q(CNT3[2]), .QN(n104) );
  DFFRX2 \CNT3_reg[1]  ( .D(n887), .CK(clk), .RN(n1047), .Q(CNT3[1]), .QN(n105) );
  DFFRX2 \CNT3_reg[0]  ( .D(n888), .CK(clk), .RN(n1047), .Q(CNT3[0]), .QN(n106) );
  DFFRX2 \CNT4_reg[7]  ( .D(n897), .CK(clk), .RN(n1048), .Q(CNT4[7]), .QN(n83)
         );
  DFFRX2 \CNT4_reg[6]  ( .D(n898), .CK(clk), .RN(n1048), .Q(CNT4[6]), .QN(n84)
         );
  DFFRX2 \CNT4_reg[5]  ( .D(n899), .CK(clk), .RN(n1048), .Q(CNT4[5]), .QN(n85)
         );
  DFFRX2 \CNT4_reg[4]  ( .D(n900), .CK(clk), .RN(n1048), .Q(CNT4[4]), .QN(n86)
         );
  DFFRX2 \CNT4_reg[3]  ( .D(n901), .CK(clk), .RN(n1048), .Q(CNT4[3]), .QN(n87)
         );
  DFFRX2 \CNT4_reg[2]  ( .D(n902), .CK(clk), .RN(n1048), .Q(CNT4[2]), .QN(n88)
         );
  DFFRX2 \CNT4_reg[1]  ( .D(n903), .CK(clk), .RN(n1084), .Q(CNT4[1]), .QN(n89)
         );
  DFFRX2 \CNT4_reg[0]  ( .D(n904), .CK(clk), .RN(n1084), .Q(CNT4[0]), .QN(n90)
         );
  DFFRX2 \CNT5_reg[0]  ( .D(n896), .CK(clk), .RN(n1048), .Q(CNT5[0]), .QN(n98)
         );
  DFFQX2 \HC1_reg[0]  ( .D(n636), .CK(clk), .Q(HC1[0]) );
  DFFQX2 \HC1_reg[1]  ( .D(n629), .CK(clk), .Q(HC1[1]) );
  DFFQX2 \M1_reg[7]  ( .D(n661), .CK(clk), .Q(M1[7]) );
  DFFRX2 \CNT5_reg[7]  ( .D(n889), .CK(clk), .RN(n1047), .Q(CNT5[7]), .QN(n91)
         );
  DFFRX2 \CNT5_reg[4]  ( .D(n892), .CK(clk), .RN(n1048), .Q(CNT5[4]), .QN(n94)
         );
  DFFRX2 \CNT5_reg[5]  ( .D(n891), .CK(clk), .RN(n1048), .Q(CNT5[5]), .QN(n93)
         );
  DFFRX2 \CNT5_reg[6]  ( .D(n890), .CK(clk), .RN(n1047), .Q(CNT5[6]), .QN(n92)
         );
  DFFQX1 \tmp_T0_reg[1]  ( .D(n721), .CK(clk), .Q(tmp_T0[1]) );
  DFFQX1 \tmp_T0_reg[3]  ( .D(n713), .CK(clk), .Q(tmp_T0[3]) );
  DFFQX1 \tmp_T0_reg[2]  ( .D(n717), .CK(clk), .Q(tmp_T0[2]) );
  DFFQX1 \tmp_T0_reg[0]  ( .D(n725), .CK(clk), .Q(tmp_T0[0]) );
  DFFQX1 \tmp_T1_reg[3]  ( .D(n729), .CK(clk), .Q(tmp_T1[3]) );
  DFFQX1 \tmp_T1_reg[1]  ( .D(n737), .CK(clk), .Q(tmp_T1[1]) );
  DFFQX1 \tmp_T1_reg[2]  ( .D(n733), .CK(clk), .Q(tmp_T1[2]) );
  DFFQX1 \tmp_T1_reg[0]  ( .D(n741), .CK(clk), .Q(tmp_T1[0]) );
  DFFQX1 \node_reg[2]  ( .D(n646), .CK(clk), .Q(node[2]) );
  DFFQX1 \node_reg[1]  ( .D(n647), .CK(clk), .Q(node[1]) );
  DFFQX1 \node_reg[0]  ( .D(n648), .CK(clk), .Q(node[0]) );
  DFFX1 \node_reg[3]  ( .D(n645), .CK(clk), .QN(n277) );
  DFFRX1 \cnt_reg[6]  ( .D(n857), .CK(clk), .RN(n1045), .Q(cnt[6]) );
  DFFQX1 \RegB_v_reg[7]  ( .D(n842), .CK(clk), .Q(RegB_v[7]) );
  DFFRX1 \cnt_reg[3]  ( .D(n846), .CK(clk), .RN(n1046), .Q(cnt[3]) );
  DFFRX1 \cnt_reg[4]  ( .D(n845), .CK(clk), .RN(n1046), .Q(cnt[4]) );
  DFFRX1 \cnt_reg[5]  ( .D(n844), .CK(clk), .RN(n1046), .Q(cnt[5]) );
  DFFRX2 \CNT5_reg[1]  ( .D(n895), .CK(clk), .RN(n1048), .Q(CNT5[1]), .QN(n97)
         );
  DFFRX2 \int_j_reg[0]  ( .D(n850), .CK(clk), .RN(n1045), .Q(int_j[0]), .QN(
        n252) );
  DFFRX2 \CNT5_reg[2]  ( .D(n894), .CK(clk), .RN(n1048), .Q(CNT5[2]), .QN(n96)
         );
  DFFRX2 \CNT5_reg[3]  ( .D(n893), .CK(clk), .RN(n1048), .Q(CNT5[3]), .QN(n95)
         );
  DFFRX1 \cnt2_reg[1]  ( .D(n853), .CK(clk), .RN(n1046), .Q(cnt2[1]), .QN(n150) );
  DFFRX1 \cnt2_reg[0]  ( .D(n852), .CK(clk), .RN(n1046), .Q(cnt2[0]), .QN(n151) );
  DFFQX1 \RegA_t_reg[2]  ( .D(n774), .CK(clk), .Q(RegA_t[2]) );
  DFFX1 \tmp_HC_reg[3]  ( .D(n616), .CK(clk), .Q(tmp_HC[3]), .QN(n285) );
  DFFX1 \tmp_HC_reg[4]  ( .D(n609), .CK(clk), .Q(tmp_HC[4]), .QN(n284) );
  DFFX1 \tmp_HC_reg[5]  ( .D(n602), .CK(clk), .Q(tmp_HC[5]), .QN(n283) );
  DFFX1 \tmp_HC_reg[6]  ( .D(n595), .CK(clk), .Q(tmp_HC[6]), .QN(n282) );
  DFFX1 \tmp_HC_reg[7]  ( .D(n644), .CK(clk), .Q(tmp_HC[7]), .QN(n281) );
  DFFX1 \tmp_MK_reg[7]  ( .D(n662), .CK(clk), .Q(n1017), .QN(n289) );
  DFFX1 \tmp_HC_reg[1]  ( .D(n630), .CK(clk), .Q(tmp_HC[1]), .QN(n287) );
  DFFX1 \tmp_HC_reg[2]  ( .D(n623), .CK(clk), .Q(tmp_HC[2]), .QN(n286) );
  DFFX1 \tmp_HC_reg[0]  ( .D(n637), .CK(clk), .Q(tmp_HC[0]), .QN(n288) );
  DFFQX1 \RegA_v_reg[4]  ( .D(n836), .CK(clk), .Q(RegA_v[4]) );
  DFFQX1 \RegA_v_reg[5]  ( .D(n835), .CK(clk), .Q(RegA_v[5]) );
  DFFQX1 \RegA_v_reg[6]  ( .D(n834), .CK(clk), .Q(RegA_v[6]) );
  DFFQX1 \RegA_v_reg[2]  ( .D(n838), .CK(clk), .Q(RegA_v[2]) );
  DFFRX2 \CNT1_reg[7]  ( .D(n865), .CK(clk), .RN(n1084), .Q(CNT1[7]), .QN(n115) );
  DFFRX2 \CNT2_reg[7]  ( .D(n905), .CK(clk), .RN(n1084), .Q(CNT2[7]), .QN(n75)
         );
  DFFRX2 \CNT1_reg[6]  ( .D(n866), .CK(clk), .RN(n1084), .Q(CNT1[6]), .QN(n116) );
  DFFRX2 \CNT1_reg[5]  ( .D(n867), .CK(clk), .RN(n1084), .Q(CNT1[5]), .QN(n117) );
  DFFRX2 \CNT1_reg[4]  ( .D(n868), .CK(clk), .RN(n1084), .Q(CNT1[4]), .QN(n118) );
  DFFRX2 \CNT1_reg[3]  ( .D(n869), .CK(clk), .RN(n1084), .Q(CNT1[3]), .QN(n119) );
  DFFRX2 \CNT2_reg[6]  ( .D(n906), .CK(clk), .RN(n1084), .Q(CNT2[6]), .QN(n76)
         );
  DFFRX2 \CNT2_reg[5]  ( .D(n907), .CK(clk), .RN(n1084), .Q(CNT2[5]), .QN(n77)
         );
  DFFRX2 \CNT2_reg[4]  ( .D(n908), .CK(clk), .RN(n1084), .Q(CNT2[4]), .QN(n78)
         );
  DFFRX2 \CNT2_reg[3]  ( .D(n909), .CK(clk), .RN(n1084), .Q(CNT2[3]), .QN(n79)
         );
  DFFRX2 \CNT1_reg[2]  ( .D(n870), .CK(clk), .RN(n1084), .Q(CNT1[2]), .QN(n120) );
  DFFRX2 \CNT1_reg[1]  ( .D(n871), .CK(clk), .RN(n1084), .Q(CNT1[1]), .QN(n121) );
  DFFRX2 \CNT2_reg[2]  ( .D(n910), .CK(clk), .RN(n1084), .Q(CNT2[2]), .QN(n80)
         );
  DFFRX2 \CNT2_reg[1]  ( .D(n911), .CK(clk), .RN(n1084), .Q(CNT2[1]), .QN(n81)
         );
  DFFRX2 \CNT1_reg[0]  ( .D(n872), .CK(clk), .RN(n1084), .Q(CNT1[0]), .QN(n122) );
  DFFRX2 \CNT2_reg[0]  ( .D(n912), .CK(clk), .RN(n1084), .Q(CNT2[0]), .QN(n82)
         );
  DFFQX1 \RegB_v_reg[5]  ( .D(n782), .CK(clk), .Q(RegB_v[5]) );
  EDFFXL \Tree_0_reg[0][1]  ( .D(n1112), .E(n1023), .CK(clk), .QN(n271) );
  EDFFXL \Tree_1_reg[0][1]  ( .D(n1114), .E(n1023), .CK(clk), .QN(n263) );
  EDFFXL \Tree_0_reg[0][3]  ( .D(n1119), .E(n1023), .CK(clk), .QN(n269) );
  EDFFXL \Tree_1_reg[0][3]  ( .D(n1116), .E(n1023), .CK(clk), .QN(n261) );
  EDFFXL \Tree_0_reg[0][2]  ( .D(n1118), .E(n1023), .CK(clk), .QN(n270) );
  EDFFXL \Tree_1_reg[0][2]  ( .D(n1115), .E(n1023), .CK(clk), .QN(n262) );
  EDFFXL \Tree_0_reg[0][0]  ( .D(n1117), .E(n1023), .CK(clk), .QN(n272) );
  EDFFXL \Tree_1_reg[0][0]  ( .D(n1113), .E(n1023), .CK(clk), .QN(n264) );
  EDFFXL \Tree_0_reg[3][1]  ( .D(n1112), .E(n1024), .CK(clk), .QN(n275) );
  EDFFXL \Tree_1_reg[3][1]  ( .D(n1114), .E(n1024), .CK(clk), .QN(n267) );
  EDFFXL \Tree_0_reg[3][3]  ( .D(n1119), .E(n1024), .CK(clk), .QN(n273) );
  EDFFXL \Tree_1_reg[3][3]  ( .D(n1116), .E(n1024), .CK(clk), .QN(n265) );
  EDFFXL \Tree_0_reg[3][2]  ( .D(n1118), .E(n1024), .CK(clk), .QN(n274) );
  EDFFXL \Tree_1_reg[3][2]  ( .D(n1115), .E(n1024), .CK(clk), .QN(n266) );
  EDFFXL \Tree_0_reg[3][0]  ( .D(n1117), .E(n1024), .CK(clk), .QN(n276) );
  EDFFXL \Tree_1_reg[3][0]  ( .D(n1113), .E(n1024), .CK(clk), .QN(n268) );
  DFFXL \addnum_reg[7]  ( .D(n649), .CK(clk), .Q(addnum[7]), .QN(n297) );
  DFFQXL \ListB_reg[3][1]  ( .D(n816), .CK(clk), .Q(\ListB[3][1] ) );
  DFFQXL \ListB_reg[3][2]  ( .D(n815), .CK(clk), .Q(\ListB[3][2] ) );
  DFFQXL \ListB_reg[3][3]  ( .D(n814), .CK(clk), .Q(\ListB[3][3] ) );
  DFFQXL \ListB_reg[3][4]  ( .D(n813), .CK(clk), .Q(\ListB[3][4] ) );
  DFFQXL \ListB_reg[3][5]  ( .D(n812), .CK(clk), .Q(\ListB[3][5] ) );
  DFFQXL \ListB_reg[3][6]  ( .D(n811), .CK(clk), .Q(\ListB[3][6] ) );
  DFFQXL \ListA_reg[5][1]  ( .D(n771), .CK(clk), .Q(\ListA[5][1] ) );
  DFFQXL \ListA_reg[2][1]  ( .D(n759), .CK(clk), .Q(\ListA[2][1] ) );
  DFFQXL \ListA_reg[2][2]  ( .D(n758), .CK(clk), .Q(\ListA[2][2] ) );
  DFFQXL \ListA_reg[5][2]  ( .D(n770), .CK(clk), .Q(\ListA[5][2] ) );
  DFFQXL \ListA_reg[2][0]  ( .D(n760), .CK(clk), .Q(\ListA[2][0] ) );
  DFFQXL \ListA_reg[5][0]  ( .D(n772), .CK(clk), .Q(\ListA[5][0] ) );
  DFFQXL \ListB_reg[2][7]  ( .D(n802), .CK(clk), .Q(\ListB[2][7] ) );
  DFFQXL \ListB_reg[2][0]  ( .D(n809), .CK(clk), .Q(\ListB[2][0] ) );
  DFFQXL \ListB_reg[5][0]  ( .D(n833), .CK(clk), .Q(\ListB[5][0] ) );
  DFFQXL \ListB_reg[2][1]  ( .D(n808), .CK(clk), .Q(\ListB[2][1] ) );
  DFFQXL \ListB_reg[5][1]  ( .D(n832), .CK(clk), .Q(\ListB[5][1] ) );
  DFFQXL \ListB_reg[2][2]  ( .D(n807), .CK(clk), .Q(\ListB[2][2] ) );
  DFFQXL \ListB_reg[5][2]  ( .D(n831), .CK(clk), .Q(\ListB[5][2] ) );
  DFFQXL \ListB_reg[2][3]  ( .D(n806), .CK(clk), .Q(\ListB[2][3] ) );
  DFFQXL \ListB_reg[5][3]  ( .D(n830), .CK(clk), .Q(\ListB[5][3] ) );
  DFFQXL \ListB_reg[2][4]  ( .D(n805), .CK(clk), .Q(\ListB[2][4] ) );
  DFFQXL \ListB_reg[5][4]  ( .D(n829), .CK(clk), .Q(\ListB[5][4] ) );
  DFFQXL \ListB_reg[2][5]  ( .D(n804), .CK(clk), .Q(\ListB[2][5] ) );
  DFFQXL \ListB_reg[5][5]  ( .D(n828), .CK(clk), .Q(\ListB[5][5] ) );
  DFFQXL \ListB_reg[2][6]  ( .D(n803), .CK(clk), .Q(\ListB[2][6] ) );
  DFFQXL \ListB_reg[5][7]  ( .D(n826), .CK(clk), .Q(\ListB[5][7] ) );
  DFFQXL \ListB_reg[5][6]  ( .D(n827), .CK(clk), .Q(\ListB[5][6] ) );
  DFFQXL \ListB_reg[1][1]  ( .D(n800), .CK(clk), .Q(\ListB[1][1] ) );
  DFFQXL \ListB_reg[1][2]  ( .D(n799), .CK(clk), .Q(\ListB[1][2] ) );
  DFFQXL \ListB_reg[1][3]  ( .D(n798), .CK(clk), .Q(\ListB[1][3] ) );
  DFFQXL \ListB_reg[1][4]  ( .D(n797), .CK(clk), .Q(\ListB[1][4] ) );
  DFFQXL \ListB_reg[1][5]  ( .D(n796), .CK(clk), .Q(\ListB[1][5] ) );
  DFFQXL \ListB_reg[1][6]  ( .D(n795), .CK(clk), .Q(\ListB[1][6] ) );
  DFFXL \addnum_reg[5]  ( .D(n651), .CK(clk), .Q(addnum[5]), .QN(n299) );
  DFFXL \addnum_reg[6]  ( .D(n650), .CK(clk), .Q(addnum[6]), .QN(n298) );
  DFFQXL \ListA_reg[3][1]  ( .D(n763), .CK(clk), .Q(\ListA[3][1] ) );
  DFFQXL \ListA_reg[0][1]  ( .D(n750), .CK(clk), .Q(\ListA[0][1] ) );
  DFFQXL \ListA_reg[0][3]  ( .D(n746), .CK(clk), .Q(\ListA[0][3] ) );
  DFFQXL \ListA_reg[3][3]  ( .D(n761), .CK(clk), .Q(\ListA[3][3] ) );
  DFFQXL \ListA_reg[0][2]  ( .D(n748), .CK(clk), .Q(\ListA[0][2] ) );
  DFFQXL \ListA_reg[3][2]  ( .D(n762), .CK(clk), .Q(\ListA[3][2] ) );
  DFFQXL \ListA_reg[0][0]  ( .D(n752), .CK(clk), .Q(\ListA[0][0] ) );
  DFFQXL \ListA_reg[3][0]  ( .D(n764), .CK(clk), .Q(\ListA[3][0] ) );
  DFFQXL \ListB_reg[3][7]  ( .D(n810), .CK(clk), .Q(\ListB[3][7] ) );
  DFFQXL \ListB_reg[3][0]  ( .D(n817), .CK(clk), .Q(\ListB[3][0] ) );
  DFFQXL \ListA_reg[2][3]  ( .D(n757), .CK(clk), .Q(\ListA[2][3] ) );
  DFFQXL \ListA_reg[5][3]  ( .D(n769), .CK(clk), .Q(\ListA[5][3] ) );
  DFFQXL \ListA_reg[1][1]  ( .D(n755), .CK(clk), .Q(\ListA[1][1] ) );
  DFFQXL \ListA_reg[1][3]  ( .D(n753), .CK(clk), .Q(\ListA[1][3] ) );
  DFFQXL \ListA_reg[1][2]  ( .D(n754), .CK(clk), .Q(\ListA[1][2] ) );
  DFFQXL \ListA_reg[1][0]  ( .D(n756), .CK(clk), .Q(\ListA[1][0] ) );
  DFFQXL \ListB_reg[4][7]  ( .D(n818), .CK(clk), .Q(\ListB[4][7] ) );
  DFFQXL \ListB_reg[1][0]  ( .D(n801), .CK(clk), .Q(\ListB[1][0] ) );
  DFFQXL \ListB_reg[1][7]  ( .D(n794), .CK(clk), .Q(\ListB[1][7] ) );
  DFFXL \addnum_reg[3]  ( .D(n653), .CK(clk), .Q(addnum[3]), .QN(n301) );
  DFFXL \addnum_reg[4]  ( .D(n652), .CK(clk), .Q(addnum[4]), .QN(n300) );
  DFFXL \addnum_reg[1]  ( .D(n655), .CK(clk), .Q(addnum[1]), .QN(n303) );
  DFFXL \addnum_reg[2]  ( .D(n654), .CK(clk), .Q(addnum[2]), .QN(n302) );
  DFFXL \addnum_reg[0]  ( .D(n705), .CK(clk), .Q(addnum[0]), .QN(n304) );
  DFFQX1 \RegA_v_reg[7]  ( .D(n841), .CK(clk), .Q(RegA_v[7]) );
  DFFRX1 \int_j_reg[1]  ( .D(n849), .CK(clk), .RN(n1046), .Q(int_j[1]), .QN(
        n251) );
  DFFRX1 \int_i_reg[1]  ( .D(n847), .CK(clk), .RN(n1046), .Q(int_i[1]), .QN(
        n259) );
  DFFRX1 \int_j_reg[2]  ( .D(n858), .CK(clk), .RN(n1045), .Q(int_j[2]), .QN(
        n249) );
  DFFRX1 \int_k_reg[2]  ( .D(n859), .CK(clk), .RN(n1046), .Q(\int_k[2] ), .QN(
        n253) );
  DFFRX1 \int_i_reg[0]  ( .D(n848), .CK(clk), .RN(n1046), .Q(int_i[0]), .QN(
        n260) );
  DFFRX1 \cnt_reg[2]  ( .D(n854), .CK(clk), .RN(n1046), .Q(cnt[2]), .QN(n139)
         );
  DFFRX1 \int_k_reg[0]  ( .D(n861), .CK(clk), .RN(n1045), .Q(N488), .QN(n256)
         );
  DFFQX1 \RegA_v_reg[3]  ( .D(n837), .CK(clk), .Q(RegA_v[3]) );
  DFFRX1 \cnt_reg[0]  ( .D(n856), .CK(clk), .RN(n1045), .Q(cnt[0]), .QN(n149)
         );
  DFFQX1 \RegB_v_reg[4]  ( .D(n784), .CK(clk), .Q(RegB_v[4]) );
  DFFQX1 \RegB_t_reg[3]  ( .D(n745), .CK(clk), .Q(RegB_t[3]) );
  DFFQX1 \RegB_v_reg[2]  ( .D(n788), .CK(clk), .Q(RegB_v[2]) );
  DFFRX4 \cs_reg[1]  ( .D(n863), .CK(clk), .RN(n1045), .Q(cs[1]), .QN(n310) );
  DFFRX4 \cs_reg[2]  ( .D(n862), .CK(clk), .RN(n1045), .Q(cs[2]), .QN(n309) );
  DFFRX1 \int_i_reg[2]  ( .D(n851), .CK(clk), .RN(n1046), .Q(int_i[2]), .QN(
        n258) );
  DFFX1 \L_idx_reg[0]  ( .D(n779), .CK(clk), .QN(n248) );
  DFFX1 \L_idx_reg[1]  ( .D(n778), .CK(clk), .QN(n247) );
  DFFX1 \L_idx_reg[2]  ( .D(n777), .CK(clk), .QN(n246) );
  DFFQXL \ListA_reg[4][3]  ( .D(n765), .CK(clk), .Q(\ListA[4][3] ) );
  DFFQXL \ListA_reg[4][1]  ( .D(n767), .CK(clk), .Q(\ListA[4][1] ) );
  DFFQXL \ListA_reg[4][2]  ( .D(n766), .CK(clk), .Q(\ListA[4][2] ) );
  DFFQXL \ListA_reg[4][0]  ( .D(n768), .CK(clk), .Q(\ListA[4][0] ) );
  DFFQXL \Tree_1_reg[4][0]  ( .D(n742), .CK(clk), .Q(\Tree_1[4][0] ) );
  DFFQXL \Tree_1_reg[2][0]  ( .D(n743), .CK(clk), .Q(\Tree_1[2][0] ) );
  DFFQXL \Tree_1_reg[1][0]  ( .D(n744), .CK(clk), .Q(\Tree_1[1][0] ) );
  DFFQXL \Tree_1_reg[4][3]  ( .D(n730), .CK(clk), .Q(\Tree_1[4][3] ) );
  DFFQXL \Tree_1_reg[4][2]  ( .D(n734), .CK(clk), .Q(\Tree_1[4][2] ) );
  DFFQXL \Tree_1_reg[4][1]  ( .D(n738), .CK(clk), .Q(\Tree_1[4][1] ) );
  DFFQXL \Tree_1_reg[2][3]  ( .D(n731), .CK(clk), .Q(\Tree_1[2][3] ) );
  DFFQXL \Tree_1_reg[2][2]  ( .D(n735), .CK(clk), .Q(\Tree_1[2][2] ) );
  DFFQXL \Tree_1_reg[2][1]  ( .D(n739), .CK(clk), .Q(\Tree_1[2][1] ) );
  DFFQXL \Tree_1_reg[1][3]  ( .D(n732), .CK(clk), .Q(\Tree_1[1][3] ) );
  DFFQXL \Tree_1_reg[1][2]  ( .D(n736), .CK(clk), .Q(\Tree_1[1][2] ) );
  DFFQXL \Tree_1_reg[1][1]  ( .D(n740), .CK(clk), .Q(\Tree_1[1][1] ) );
  DFFQXL \Tree_0_reg[4][3]  ( .D(n714), .CK(clk), .Q(\Tree_0[4][3] ) );
  DFFQXL \Tree_0_reg[4][2]  ( .D(n718), .CK(clk), .Q(\Tree_0[4][2] ) );
  DFFQXL \Tree_0_reg[4][1]  ( .D(n722), .CK(clk), .Q(\Tree_0[4][1] ) );
  DFFQXL \Tree_0_reg[4][0]  ( .D(n726), .CK(clk), .Q(\Tree_0[4][0] ) );
  DFFQXL \Tree_0_reg[2][3]  ( .D(n715), .CK(clk), .Q(\Tree_0[2][3] ) );
  DFFQXL \Tree_0_reg[2][2]  ( .D(n719), .CK(clk), .Q(\Tree_0[2][2] ) );
  DFFQXL \Tree_0_reg[2][1]  ( .D(n723), .CK(clk), .Q(\Tree_0[2][1] ) );
  DFFQXL \Tree_0_reg[2][0]  ( .D(n727), .CK(clk), .Q(\Tree_0[2][0] ) );
  DFFQXL \Tree_0_reg[1][3]  ( .D(n716), .CK(clk), .Q(\Tree_0[1][3] ) );
  DFFQXL \Tree_0_reg[1][2]  ( .D(n720), .CK(clk), .Q(\Tree_0[1][2] ) );
  DFFQXL \Tree_0_reg[1][1]  ( .D(n724), .CK(clk), .Q(\Tree_0[1][1] ) );
  DFFQXL \Tree_0_reg[1][0]  ( .D(n728), .CK(clk), .Q(\Tree_0[1][0] ) );
  DFFQXL \ListB_reg[4][5]  ( .D(n820), .CK(clk), .Q(\ListB[4][5] ) );
  DFFQXL \ListB_reg[4][4]  ( .D(n821), .CK(clk), .Q(\ListB[4][4] ) );
  DFFQXL \ListB_reg[4][3]  ( .D(n822), .CK(clk), .Q(\ListB[4][3] ) );
  DFFQXL \ListB_reg[4][2]  ( .D(n823), .CK(clk), .Q(\ListB[4][2] ) );
  DFFQXL \ListB_reg[4][1]  ( .D(n824), .CK(clk), .Q(\ListB[4][1] ) );
  DFFQXL \ListB_reg[4][0]  ( .D(n825), .CK(clk), .Q(\ListB[4][0] ) );
  DFFQXL \ListB_reg[4][6]  ( .D(n819), .CK(clk), .Q(\ListB[4][6] ) );
  DFFQX2 \HC6_reg[1]  ( .D(n624), .CK(clk), .Q(HC6[1]) );
  DFFQX2 \HC6_reg[0]  ( .D(n631), .CK(clk), .Q(HC6[0]) );
  DFFQX2 \M6_reg[7]  ( .D(n656), .CK(clk), .Q(M6[7]) );
  DFFQX2 \HC3_reg[7]  ( .D(n641), .CK(clk), .Q(HC3[7]) );
  DFFQX2 \HC3_reg[4]  ( .D(n606), .CK(clk), .Q(HC3[4]) );
  DFFQX2 \HC3_reg[3]  ( .D(n613), .CK(clk), .Q(HC3[3]) );
  DFFQX2 \HC3_reg[2]  ( .D(n620), .CK(clk), .Q(HC3[2]) );
  DFFQX2 \HC3_reg[1]  ( .D(n627), .CK(clk), .Q(HC3[1]) );
  DFFQX2 \HC3_reg[0]  ( .D(n634), .CK(clk), .Q(HC3[0]) );
  DFFQX2 \M3_reg[7]  ( .D(n659), .CK(clk), .Q(M3[7]) );
  DFFQX2 \HC4_reg[7]  ( .D(n640), .CK(clk), .Q(HC4[7]) );
  DFFQX2 \HC4_reg[4]  ( .D(n605), .CK(clk), .Q(HC4[4]) );
  DFFQX2 \HC4_reg[3]  ( .D(n612), .CK(clk), .Q(HC4[3]) );
  DFFQX2 \HC4_reg[2]  ( .D(n619), .CK(clk), .Q(HC4[2]) );
  DFFQX2 \HC4_reg[1]  ( .D(n626), .CK(clk), .Q(HC4[1]) );
  DFFQX2 \HC4_reg[0]  ( .D(n633), .CK(clk), .Q(HC4[0]) );
  DFFQX2 \M4_reg[7]  ( .D(n658), .CK(clk), .Q(M4[7]) );
  DFFQX2 \HC5_reg[7]  ( .D(n639), .CK(clk), .Q(HC5[7]) );
  DFFQX2 \HC5_reg[4]  ( .D(n604), .CK(clk), .Q(HC5[4]) );
  DFFQX2 \HC5_reg[3]  ( .D(n611), .CK(clk), .Q(HC5[3]) );
  DFFQX2 \HC5_reg[2]  ( .D(n618), .CK(clk), .Q(HC5[2]) );
  DFFQX2 \HC5_reg[1]  ( .D(n625), .CK(clk), .Q(HC5[1]) );
  DFFQX2 \HC5_reg[0]  ( .D(n632), .CK(clk), .Q(HC5[0]) );
  DFFQX2 \M5_reg[7]  ( .D(n657), .CK(clk), .Q(M5[7]) );
  DFFQX2 \HC1_reg[7]  ( .D(n643), .CK(clk), .Q(HC1[7]) );
  DFFQX2 \HC1_reg[4]  ( .D(n608), .CK(clk), .Q(HC1[4]) );
  DFFQX2 \HC1_reg[3]  ( .D(n615), .CK(clk), .Q(HC1[3]) );
  DFFQX2 \HC1_reg[2]  ( .D(n622), .CK(clk), .Q(HC1[2]) );
  DFFRX2 CNT_valid_reg ( .D(N774), .CK(clk), .RN(n1084), .Q(CNT_valid) );
  DFFQX1 \RegB_v_reg[6]  ( .D(n780), .CK(clk), .Q(RegB_v[6]) );
  DFFQX1 \RegB_v_reg[3]  ( .D(n786), .CK(clk), .Q(RegB_v[3]) );
  DFFRX2 \cs_reg[0]  ( .D(n864), .CK(clk), .RN(n1045), .Q(cs[0]), .QN(n311) );
  DFFQX1 \RegA_v_reg[1]  ( .D(n839), .CK(clk), .Q(RegA_v[1]) );
  DFFQX1 \RegA_v_reg[0]  ( .D(n840), .CK(clk), .Q(RegA_v[0]) );
  DFFQX1 \RegB_v_reg[1]  ( .D(n790), .CK(clk), .Q(RegB_v[1]) );
  DFFQX1 \RegB_v_reg[0]  ( .D(n792), .CK(clk), .Q(RegB_v[0]) );
  DFFRX2 \cnt_reg[1]  ( .D(n855), .CK(clk), .RN(n1045), .Q(cnt[1]), .QN(n140)
         );
  DFFQX2 \RegA_t_reg[1]  ( .D(n775), .CK(clk), .Q(RegA_t[1]) );
  DFFQX2 \RegB_t_reg[1]  ( .D(n749), .CK(clk), .Q(RegB_t[1]) );
  DFFQX2 \RegB_t_reg[0]  ( .D(n751), .CK(clk), .Q(RegB_t[0]) );
  DFFQX2 \RegB_t_reg[2]  ( .D(n747), .CK(clk), .Q(RegB_t[2]) );
  INVX1 U745 ( .A(net7476), .Y(n914) );
  INVX6 U746 ( .A(net7492), .Y(net7476) );
  OAI21X2 U748 ( .A0(RegA_v[6]), .A1(n1213), .B0(n493), .Y(n492) );
  NAND2X4 U749 ( .A(n952), .B(n502), .Y(n501) );
  NOR2X1 U750 ( .A(n451), .B(n916), .Y(n960) );
  NAND2X6 U751 ( .A(n1037), .B(n422), .Y(n916) );
  OAI21X2 U752 ( .A0(RegB_v[7]), .A1(n1153), .B0(n490), .Y(n360) );
  INVX3 U753 ( .A(RegB_t[1]), .Y(n1120) );
  NAND2X4 U754 ( .A(gray_data[2]), .B(gray_data[1]), .Y(net5501) );
  NOR2X4 U755 ( .A(gray_data[0]), .B(gray_data[2]), .Y(n938) );
  NAND2X6 U756 ( .A(net5452), .B(net7189), .Y(n915) );
  INVX1 U760 ( .A(RegA_v[0]), .Y(n1168) );
  CLKINVX1 U762 ( .A(n388), .Y(n1104) );
  NOR2X2 U763 ( .A(n980), .B(N488), .Y(n388) );
  INVX1 U764 ( .A(RegB_t[0]), .Y(n1149) );
  INVX3 U765 ( .A(RegA_t[2]), .Y(n1134) );
  OAI2BB2X1 U766 ( .B0(n569), .B1(n574), .A0N(n569), .A1N(cs[0]), .Y(n864) );
  CLKINVX1 U767 ( .A(n457), .Y(n1102) );
  OAI221X4 U768 ( .A0(n251), .A1(n523), .B0(n996), .B1(n247), .C0(n524), .Y(
        n457) );
  OAI21X4 U769 ( .A0(RegA_t[2]), .A1(n1141), .B0(n508), .Y(n507) );
  NAND2X2 U770 ( .A(n955), .B(n509), .Y(n508) );
  NAND2X6 U771 ( .A(cnt[1]), .B(n1044), .Y(n543) );
  NAND2X4 U772 ( .A(n957), .B(n943), .Y(n497) );
  NAND2X2 U773 ( .A(n942), .B(n500), .Y(n944) );
  CLKINVX1 U774 ( .A(n514), .Y(n1093) );
  CLKINVX1 U775 ( .A(n543), .Y(n939) );
  NOR3X4 U776 ( .A(n311), .B(cs[2]), .C(n310), .Y(n526) );
  CLKBUFX3 U777 ( .A(n429), .Y(n1035) );
  BUFX12 U778 ( .A(cnt[0]), .Y(n1044) );
  NAND2X1 U779 ( .A(n1110), .B(n999), .Y(n524) );
  BUFX4 U780 ( .A(n1100), .Y(n1031) );
  NAND2X2 U781 ( .A(n1031), .B(n455), .Y(n982) );
  NAND2X6 U782 ( .A(n1041), .B(n455), .Y(n984) );
  NAND2X6 U783 ( .A(n1010), .B(n1041), .Y(n994) );
  NAND2X6 U784 ( .A(n1010), .B(n1040), .Y(n992) );
  NAND2X6 U785 ( .A(n1040), .B(n455), .Y(n983) );
  NAND2X6 U786 ( .A(n1039), .B(n455), .Y(n981) );
  NAND2X6 U787 ( .A(n1010), .B(n1039), .Y(n993) );
  NAND2X1 U788 ( .A(n953), .B(n954), .Y(n509) );
  CLKAND2X3 U789 ( .A(n505), .B(n506), .Y(n950) );
  NAND2X1 U790 ( .A(RegB_t[3]), .B(n1127), .Y(n505) );
  NAND2X2 U791 ( .A(n948), .B(n507), .Y(n506) );
  OR2X1 U792 ( .A(RegB_t[2]), .B(n1134), .Y(n948) );
  AND2X2 U793 ( .A(RegA_t[3]), .B(n1133), .Y(n951) );
  NAND2X1 U794 ( .A(n958), .B(n501), .Y(n500) );
  NAND2X1 U795 ( .A(n1184), .B(RegB_v[2]), .Y(n958) );
  OR2X1 U796 ( .A(RegB_v[2]), .B(n1184), .Y(n942) );
  NAND2X2 U797 ( .A(n947), .B(n496), .Y(n495) );
  OR2X1 U798 ( .A(RegB_v[4]), .B(n962), .Y(n947) );
  NAND2X2 U799 ( .A(n963), .B(n497), .Y(n496) );
  OR2X1 U800 ( .A(RegA_v[5]), .B(n1205), .Y(n945) );
  INVX4 U801 ( .A(net7390), .Y(net7595) );
  OAI21X2 U802 ( .A0(RegA_v[7]), .A1(n1160), .B0(n491), .Y(n490) );
  OR2X4 U803 ( .A(n543), .B(n522), .Y(n980) );
  NAND2X1 U804 ( .A(n521), .B(n151), .Y(n517) );
  CLKBUFX3 U805 ( .A(n355), .Y(n1042) );
  AOI32X1 U806 ( .A0(n1102), .A1(n461), .A2(n1101), .B0(n462), .B1(n1010), .Y(
        n413) );
  AND2X2 U808 ( .A(n484), .B(n485), .Y(n451) );
  NAND2X1 U809 ( .A(n541), .B(n542), .Y(n531) );
  OA21XL U810 ( .A0(n1088), .A1(n252), .B0(n537), .Y(n534) );
  NAND2X2 U811 ( .A(n1010), .B(n1038), .Y(n998) );
  NAND2X2 U813 ( .A(n1010), .B(n1032), .Y(n995) );
  NOR2BX2 U814 ( .AN(n1043), .B(n1050), .Y(n320) );
  CLKINVX1 U815 ( .A(RegB_t[2]), .Y(n1141) );
  CLKINVX1 U816 ( .A(RegA_t[1]), .Y(n1121) );
  INVX3 U817 ( .A(n548), .Y(n1085) );
  OAI31XL U818 ( .A0(n549), .A1(n1010), .A2(n550), .B0(n1086), .Y(n548) );
  CLKINVX12 U819 ( .A(n934), .Y(net7156) );
  NAND2X1 U820 ( .A(n919), .B(n1012), .Y(n776) );
  OAI222XL U821 ( .A0(n453), .A1(n984), .B0(n994), .B1(n75), .C0(n1041), .C1(
        n1154), .Y(n794) );
  OAI222XL U822 ( .A0(n453), .A1(n982), .B0(n918), .B1(n91), .C0(n1031), .C1(
        n1157), .Y(n818) );
  OAI222XL U823 ( .A0(n453), .A1(n981), .B0(n993), .B1(n83), .C0(n1039), .C1(
        n1156), .Y(n810) );
  OAI222XL U824 ( .A0(n453), .A1(n983), .B0(n992), .B1(n99), .C0(n1040), .C1(
        n1155), .Y(n802) );
  CLKINVX1 U825 ( .A(n385), .Y(n1113) );
  CLKINVX1 U826 ( .A(n369), .Y(n1117) );
  CLKINVX1 U827 ( .A(n375), .Y(n1115) );
  CLKINVX1 U828 ( .A(n363), .Y(n1118) );
  CLKINVX1 U829 ( .A(n372), .Y(n1116) );
  CLKINVX1 U830 ( .A(n354), .Y(n1119) );
  CLKINVX1 U831 ( .A(n378), .Y(n1114) );
  CLKINVX1 U832 ( .A(n366), .Y(n1112) );
  CLKINVX4 U833 ( .A(reset), .Y(n1084) );
  OR2X1 U834 ( .A(cs[0]), .B(n310), .Y(n917) );
  NAND2X2 U835 ( .A(n1010), .B(n1031), .Y(n918) );
  AND2X2 U836 ( .A(n1011), .B(n1013), .Y(n919) );
  CLKINVX1 U837 ( .A(RegB_v[3]), .Y(n956) );
  CLKMX2X4 U838 ( .A(CNT5[6]), .B(N416), .S0(net5661), .Y(n890) );
  CLKMX2X4 U839 ( .A(CNT5[5]), .B(N415), .S0(net5661), .Y(n891) );
  CLKMX2X4 U840 ( .A(CNT5[4]), .B(N414), .S0(net5661), .Y(n892) );
  CLKMX2X4 U841 ( .A(CNT5[7]), .B(N417), .S0(net5661), .Y(n889) );
  BUFX16 U842 ( .A(gray_data[1]), .Y(net7390) );
  CLKMX2X4 U843 ( .A(CNT5[0]), .B(N410), .S0(net5661), .Y(n896) );
  OAI21X2 U844 ( .A0(RegB_v[6]), .A1(n1214), .B0(n492), .Y(n491) );
  NAND3X1 U845 ( .A(n383), .B(n139), .C(n526), .Y(n488) );
  NAND2X8 U862 ( .A(net7189), .B(net5500), .Y(n940) );
  MXI2X2 U863 ( .A(n114), .B(n1073), .S0(n1009), .Y(n880) );
  NOR2X8 U864 ( .A(net7595), .B(n935), .Y(net5452) );
  CLKINVX12 U866 ( .A(n941), .Y(net5661) );
  INVX1 U869 ( .A(N387), .Y(n1082) );
  INVX1 U870 ( .A(N388), .Y(n1081) );
  INVX1 U871 ( .A(N389), .Y(n1080) );
  INVX1 U872 ( .A(N390), .Y(n1079) );
  INVX1 U873 ( .A(N391), .Y(n1078) );
  INVX1 U874 ( .A(N392), .Y(n1077) );
  INVX1 U875 ( .A(N393), .Y(n1076) );
  NAND2X4 U877 ( .A(net7492), .B(gray_data[2]), .Y(n937) );
  NAND2X2 U878 ( .A(gray_data[0]), .B(net7492), .Y(net7469) );
  NOR3X4 U879 ( .A(n937), .B(gray_data[1]), .C(gray_data[0]), .Y(n936) );
  AND3X2 U880 ( .A(n331), .B(n939), .C(int_i[2]), .Y(n562) );
  MXI2X4 U881 ( .A(n90), .B(n1075), .S0(net7156), .Y(n904) );
  CLKMX2X6 U882 ( .A(CNT4[6]), .B(N408), .S0(net7156), .Y(n898) );
  CLKMX2X6 U883 ( .A(CNT4[4]), .B(N406), .S0(net7156), .Y(n900) );
  CLKMX2X6 U884 ( .A(CNT4[2]), .B(N404), .S0(net7156), .Y(n902) );
  CLKMX2X6 U885 ( .A(CNT4[5]), .B(N407), .S0(net7156), .Y(n899) );
  CLKMX2X6 U886 ( .A(CNT4[3]), .B(N405), .S0(net7156), .Y(n901) );
  CLKMX2X6 U887 ( .A(CNT4[1]), .B(N403), .S0(net7156), .Y(n903) );
  CLKMX2X6 U888 ( .A(CNT4[7]), .B(N409), .S0(net7156), .Y(n897) );
  CLKINVX20 U890 ( .A(n915), .Y(n1030) );
  CLKMX2X4 U891 ( .A(CNT6[7]), .B(N425), .S0(n1009), .Y(n873) );
  CLKMX2X4 U892 ( .A(CNT6[6]), .B(N424), .S0(n1009), .Y(n874) );
  CLKMX2X4 U893 ( .A(CNT6[5]), .B(N423), .S0(n1009), .Y(n875) );
  CLKMX2X4 U894 ( .A(CNT6[4]), .B(N422), .S0(n1009), .Y(n876) );
  CLKMX2X4 U895 ( .A(CNT6[3]), .B(N421), .S0(n1009), .Y(n877) );
  CLKMX2X4 U896 ( .A(CNT6[2]), .B(N420), .S0(n1009), .Y(n878) );
  CLKMX2X4 U897 ( .A(CNT6[1]), .B(N419), .S0(n1009), .Y(n879) );
  INVX1 U901 ( .A(N379), .Y(n1070) );
  INVX1 U902 ( .A(N380), .Y(n1069) );
  INVX1 U903 ( .A(N381), .Y(n1068) );
  INVX1 U904 ( .A(N382), .Y(n1067) );
  INVX1 U905 ( .A(N383), .Y(n1066) );
  INVX1 U906 ( .A(N384), .Y(n1065) );
  INVX1 U907 ( .A(N385), .Y(n1064) );
  BUFX4 U908 ( .A(n360), .Y(n1036) );
  NAND2X2 U909 ( .A(n525), .B(n526), .Y(n523) );
  AOI2BB1X2 U910 ( .A0N(n1213), .A1N(n996), .B0(n1018), .Y(n440) );
  AO22XL U911 ( .A0(N498), .A1(n999), .B0(RegA_v[6]), .B1(n985), .Y(n1018) );
  AOI2BB1X2 U912 ( .A0N(n1198), .A1N(n996), .B0(n1020), .Y(n444) );
  AO22XL U913 ( .A0(N496), .A1(n999), .B0(RegA_v[4]), .B1(n985), .Y(n1020) );
  AOI2BB1X2 U914 ( .A0N(n1205), .A1N(n996), .B0(n1019), .Y(n442) );
  AO22XL U915 ( .A0(N497), .A1(n999), .B0(RegA_v[5]), .B1(n985), .Y(n1019) );
  AOI2BB1X2 U916 ( .A0N(n1183), .A1N(n996), .B0(n1022), .Y(n448) );
  AOI2BB1X2 U917 ( .A0N(n956), .A1N(n996), .B0(n1021), .Y(n446) );
  NOR2X4 U918 ( .A(n1095), .B(n1093), .Y(n987) );
  INVX3 U919 ( .A(n513), .Y(n1095) );
  OA21X1 U920 ( .A0(n1175), .A1(n996), .B0(n1003), .Y(n450) );
  NAND3X4 U921 ( .A(n387), .B(n255), .C(n388), .Y(n1006) );
  NOR2X4 U922 ( .A(n514), .B(n1094), .Y(n1000) );
  AOI2BB1X2 U923 ( .A0N(n1167), .A1N(n996), .B0(n1004), .Y(n452) );
  AO22X1 U924 ( .A0(N492), .A1(n999), .B0(RegA_v[0]), .B1(n985), .Y(n1004) );
  OR4X2 U925 ( .A(n1002), .B(n381), .C(n382), .D(n1008), .Y(n353) );
  NAND2X2 U926 ( .A(n383), .B(n384), .Y(n1002) );
  NAND3X4 U927 ( .A(N296), .B(n1104), .C(n387), .Y(n1007) );
  NAND2X4 U928 ( .A(n324), .B(n1050), .Y(n986) );
  OR2XL U929 ( .A(n400), .B(n916), .Y(n1012) );
  OR2XL U930 ( .A(n1142), .B(n1037), .Y(n1013) );
  OAI2BB1X4 U931 ( .A0N(n1191), .A1N(RegB_v[3]), .B0(n944), .Y(n943) );
  NAND2X8 U932 ( .A(n945), .B(n495), .Y(n494) );
  NAND2X8 U933 ( .A(n946), .B(n494), .Y(n493) );
  OR2X2 U934 ( .A(RegB_v[5]), .B(n1206), .Y(n946) );
  AO22XL U935 ( .A0(n528), .A1(cnt[1]), .B0(N441), .B1(n1085), .Y(n855) );
  NOR2X8 U936 ( .A(n1044), .B(cnt[1]), .Y(n383) );
  CLKINVX3 U937 ( .A(n980), .Y(n999) );
  NOR2X4 U938 ( .A(cs[2]), .B(n917), .Y(n1010) );
  CLKINVX1 U939 ( .A(n1010), .Y(n1106) );
  CLKAND2X3 U940 ( .A(RegB_v[0]), .B(n1168), .Y(n949) );
  NOR3X8 U941 ( .A(n949), .B(n950), .C(n951), .Y(n503) );
  CLKINVX1 U942 ( .A(RegB_t[3]), .Y(n1133) );
  OAI2BB2X4 U943 ( .B0(n503), .B1(n504), .A0N(n1176), .A1N(RegB_v[1]), .Y(n502) );
  AOI2BB1X4 U944 ( .A0N(n1160), .A1N(n996), .B0(n1005), .Y(n453) );
  OR2XL U945 ( .A(RegB_v[1]), .B(n1176), .Y(n952) );
  INVX1 U946 ( .A(n336), .Y(n1090) );
  OR2XL U947 ( .A(RegB_t[1]), .B(n1121), .Y(n955) );
  OR2X4 U948 ( .A(RegA_t[1]), .B(n1120), .Y(n953) );
  OR2X4 U949 ( .A(RegA_t[0]), .B(n1149), .Y(n954) );
  NAND2X1 U950 ( .A(n956), .B(RegA_v[3]), .Y(n957) );
  INVX1 U951 ( .A(n337), .Y(n1089) );
  INVX1 U952 ( .A(n338), .Y(n1091) );
  INVX1 U953 ( .A(n384), .Y(n1087) );
  NAND2X1 U954 ( .A(n962), .B(RegB_v[4]), .Y(n963) );
  INVXL U955 ( .A(RegA_v[1]), .Y(n1176) );
  INVXL U956 ( .A(RegB_v[1]), .Y(n1175) );
  INVX1 U957 ( .A(RegA_v[3]), .Y(n1191) );
  NOR2X6 U958 ( .A(n999), .B(n1098), .Y(n985) );
  CLKBUFX3 U959 ( .A(n313), .Y(n1062) );
  CLKBUFX3 U960 ( .A(n318), .Y(n1052) );
  CLKBUFX3 U962 ( .A(n315), .Y(n1058) );
  CLKBUFX3 U963 ( .A(n314), .Y(n1060) );
  AND2X8 U964 ( .A(n990), .B(n1036), .Y(n989) );
  INVX16 U965 ( .A(n989), .Y(n422) );
  NAND3X1 U966 ( .A(n337), .B(n1090), .C(n338), .Y(n316) );
  OA21X1 U967 ( .A0(n544), .A1(n980), .B0(n339), .Y(n324) );
  CLKBUFX3 U968 ( .A(n321), .Y(n1050) );
  AO22XL U969 ( .A0(n528), .A1(n1044), .B0(N440), .B1(n1085), .Y(n856) );
  NOR2X1 U970 ( .A(int_i[1]), .B(int_i[0]), .Y(n331) );
  INVXL U971 ( .A(RegA_v[2]), .Y(n1184) );
  NOR2XL U972 ( .A(n1167), .B(n422), .Y(n959) );
  NOR2XL U973 ( .A(n1168), .B(n1037), .Y(n961) );
  OR3X2 U974 ( .A(n959), .B(n960), .C(n961), .Y(n840) );
  INVXL U975 ( .A(RegA_v[4]), .Y(n962) );
  NAND2X4 U976 ( .A(n1099), .B(n455), .Y(n456) );
  NOR2X4 U977 ( .A(n1093), .B(n1094), .Y(n988) );
  NAND2X2 U978 ( .A(n1038), .B(n455), .Y(n997) );
  NAND2X2 U979 ( .A(n1032), .B(n455), .Y(n991) );
  BUFX12 U980 ( .A(n424), .Y(n1037) );
  OAI222XL U981 ( .A0(n1213), .A1(n422), .B0(n439), .B1(n916), .C0(n1214), 
        .C1(n1037), .Y(n834) );
  OAI222XL U982 ( .A0(n1205), .A1(n422), .B0(n441), .B1(n916), .C0(n1206), 
        .C1(n1037), .Y(n835) );
  OAI222XL U983 ( .A0(n1198), .A1(n422), .B0(n443), .B1(n916), .C0(n962), .C1(
        n1037), .Y(n836) );
  OAI222XL U984 ( .A0(n956), .A1(n422), .B0(n445), .B1(n916), .C0(n1191), .C1(
        n1037), .Y(n837) );
  OAI222XL U985 ( .A0(n1183), .A1(n422), .B0(n447), .B1(n916), .C0(n1184), 
        .C1(n1037), .Y(n838) );
  OAI222XL U986 ( .A0(n1175), .A1(n422), .B0(n449), .B1(n916), .C0(n1176), 
        .C1(n1037), .Y(n839) );
  CLKINVX1 U987 ( .A(n489), .Y(n990) );
  NAND2X8 U988 ( .A(n462), .B(n526), .Y(n996) );
  CLKBUFX2 U989 ( .A(n321), .Y(n1049) );
  NAND3X1 U990 ( .A(n311), .B(n310), .C(cs[2]), .Y(n522) );
  XNOR2X1 U991 ( .A(N488), .B(n255), .Y(n421) );
  INVX1 U992 ( .A(RegB_v[2]), .Y(n1183) );
  AOI2BB1XL U993 ( .A0N(n259), .A1N(n260), .B0(n331), .Y(n333) );
  AOI2BB1XL U994 ( .A0N(n331), .A1N(n258), .B0(n1111), .Y(n330) );
  AOI2BB2XL U995 ( .B0(n544), .B1(n567), .A0N(n1087), .A1N(n573), .Y(n571) );
  INVX1 U996 ( .A(RegB_v[6]), .Y(n1213) );
  CLKINVX1 U997 ( .A(RegB_v[7]), .Y(n1160) );
  CLKINVX1 U998 ( .A(RegA_v[5]), .Y(n1206) );
  INVX1 U999 ( .A(RegB_v[5]), .Y(n1205) );
  INVX1 U1000 ( .A(RegB_v[4]), .Y(n1198) );
  CLKINVX1 U1001 ( .A(RegA_v[6]), .Y(n1214) );
  NAND3XL U1002 ( .A(int_j[0]), .B(n562), .C(n561), .Y(n573) );
  NAND2XL U1003 ( .A(n331), .B(n258), .Y(n332) );
  XNOR2XL U1004 ( .A(int_i[0]), .B(int_j[0]), .Y(n552) );
  XNOR2XL U1005 ( .A(int_j[1]), .B(int_i[1]), .Y(n553) );
  INVXL U1006 ( .A(n560), .Y(n1088) );
  OAI211XL U1007 ( .A0(n543), .A1(n1087), .B0(n985), .C0(n555), .Y(n547) );
  AOI31XL U1008 ( .A0(n1108), .A1(n460), .A2(n551), .B0(n1097), .Y(n550) );
  NOR2XL U1010 ( .A(n980), .B(n544), .Y(n536) );
  INVXL U1011 ( .A(n525), .Y(n1108) );
  NOR2XL U1012 ( .A(n914), .B(n572), .Y(N774) );
  AND2X1 U1013 ( .A(n386), .B(n999), .Y(n387) );
  NAND3X1 U1014 ( .A(n336), .B(n1089), .C(n338), .Y(n314) );
  NAND3X1 U1015 ( .A(n336), .B(n1091), .C(n337), .Y(n313) );
  NAND3X1 U1016 ( .A(n1089), .B(n1090), .C(n338), .Y(n318) );
  NAND3X1 U1017 ( .A(n1091), .B(n1090), .C(n337), .Y(n317) );
  NAND3X1 U1018 ( .A(n1091), .B(n1089), .C(n336), .Y(n315) );
  NOR2X2 U1019 ( .A(n514), .B(n1095), .Y(n1001) );
  INVX3 U1020 ( .A(n1033), .Y(n1092) );
  NAND2XL U1021 ( .A(n577), .B(n525), .Y(n566) );
  NOR2XL U1022 ( .A(RegB_v[0]), .B(n1168), .Y(n504) );
  NOR2X4 U1023 ( .A(n139), .B(n1109), .Y(n462) );
  OAI33XL U1024 ( .A0(n456), .A1(n459), .A2(n457), .B0(n1106), .B1(cnt[2]), 
        .B2(n1109), .Y(n393) );
  OAI221X4 U1025 ( .A0(n252), .A1(n523), .B0(n996), .B1(n248), .C0(n1104), .Y(
        n459) );
  AO22XL U1026 ( .A0(n528), .A1(cnt[2]), .B0(N442), .B1(n1085), .Y(n854) );
  AO22XL U1027 ( .A0(N495), .A1(n999), .B0(RegA_v[3]), .B1(n985), .Y(n1021) );
  AO22XL U1028 ( .A0(N494), .A1(n999), .B0(RegA_v[2]), .B1(n985), .Y(n1022) );
  AOI22XL U1029 ( .A0(N493), .A1(n999), .B0(RegA_v[1]), .B1(n985), .Y(n1003)
         );
  OAI222XL U1030 ( .A0(n996), .A1(n246), .B0(n249), .B1(n523), .C0(n518), .C1(
        n980), .Y(n461) );
  AO22XL U1031 ( .A0(N499), .A1(n999), .B0(RegA_v[7]), .B1(n985), .Y(n1005) );
  NOR3XL U1032 ( .A(n980), .B(n1110), .C(n253), .Y(n420) );
  AND2X2 U1033 ( .A(n437), .B(n438), .Y(n400) );
  AND2X2 U1034 ( .A(n425), .B(n426), .Y(n392) );
  NOR2XL U1035 ( .A(N296), .B(N488), .Y(n563) );
  NOR2BXL U1036 ( .AN(n524), .B(n536), .Y(n535) );
  NOR2X1 U1037 ( .A(n259), .B(n1002), .Y(n382) );
  NOR3X1 U1038 ( .A(n311), .B(cs[1]), .C(n309), .Y(n384) );
  NOR2X1 U1039 ( .A(n260), .B(n1002), .Y(n381) );
  NOR2X1 U1040 ( .A(n252), .B(n339), .Y(n338) );
  NOR2X1 U1041 ( .A(n251), .B(n339), .Y(n337) );
  NAND2XL U1042 ( .A(n390), .B(n999), .Y(n386) );
  NOR2X1 U1043 ( .A(n249), .B(n339), .Y(n336) );
  NAND3XL U1044 ( .A(n140), .B(n139), .C(n1044), .Y(n458) );
  NAND3XL U1045 ( .A(n149), .B(n139), .C(cnt[1]), .Y(n460) );
  NAND2XL U1046 ( .A(n560), .B(n252), .Y(n533) );
  NAND3BXL U1047 ( .AN(n386), .B(n1104), .C(n255), .Y(n355) );
  NAND4XL U1048 ( .A(n1044), .B(n140), .C(cnt[2]), .D(n578), .Y(n555) );
  NAND2BXL U1049 ( .AN(n531), .B(int_i[0]), .Y(n530) );
  OAI211XL U1050 ( .A0(n256), .A1(n559), .B0(n1104), .C0(n1105), .Y(n861) );
  AOI2BB2XL U1051 ( .B0(\Tree_0[2][0] ), .B1(n352), .A0N(n353), .A1N(n272), 
        .Y(n367) );
  AOI2BB2XL U1052 ( .B0(\Tree_1[2][2] ), .B1(n352), .A0N(n353), .A1N(n262), 
        .Y(n373) );
  AOI2BB2XL U1053 ( .B0(\Tree_0[2][2] ), .B1(n352), .A0N(n353), .A1N(n270), 
        .Y(n361) );
  AOI2BB2XL U1054 ( .B0(\Tree_1[2][3] ), .B1(n352), .A0N(n353), .A1N(n261), 
        .Y(n370) );
  AOI2BB2XL U1055 ( .B0(\Tree_0[2][3] ), .B1(n352), .A0N(n353), .A1N(n269), 
        .Y(n348) );
  AOI2BB2XL U1056 ( .B0(\Tree_1[2][1] ), .B1(n352), .A0N(n353), .A1N(n263), 
        .Y(n376) );
  AOI2BB2XL U1057 ( .B0(\Tree_0[2][1] ), .B1(n352), .A0N(n353), .A1N(n271), 
        .Y(n364) );
  OAI211XL U1058 ( .A0(n252), .A1(n537), .B0(n533), .C0(n538), .Y(n850) );
  NOR2XL U1059 ( .A(n539), .B(n388), .Y(n538) );
  OAI211XL U1060 ( .A0(n310), .A1(n570), .B0(n571), .C0(n572), .Y(n568) );
  NOR2X2 U1061 ( .A(n1002), .B(n258), .Y(n1008) );
  OAI222X1 U1062 ( .A0(n249), .A1(n515), .B0(n516), .B1(n487), .C0(n258), .C1(
        n517), .Y(n513) );
  AOI2BB2XL U1063 ( .B0(\int_k[2] ), .B1(n149), .A0N(n149), .A1N(n518), .Y(
        n516) );
  OAI222X1 U1064 ( .A0(n251), .A1(n515), .B0(n519), .B1(n487), .C0(n259), .C1(
        n517), .Y(n512) );
  AOI2BB2XL U1065 ( .B0(n1044), .B1(n1110), .A0N(n255), .A1N(n1044), .Y(n519)
         );
  NAND4XL U1066 ( .A(n561), .B(n577), .C(n462), .D(int_j[0]), .Y(n564) );
  CLKBUFX3 U1067 ( .A(n391), .Y(n1033) );
  OAI211XL U1068 ( .A0(n149), .A1(n487), .B0(n515), .C0(n517), .Y(n391) );
  INVXL U1069 ( .A(RegB_v[0]), .Y(n1167) );
  OR2XL U1070 ( .A(n1149), .B(n422), .Y(n1011) );
  NOR2XL U1072 ( .A(n1133), .B(n422), .Y(n1014) );
  NOR2XL U1073 ( .A(n392), .B(n916), .Y(n1015) );
  NOR2XL U1074 ( .A(n1127), .B(n1037), .Y(n1016) );
  OR3X2 U1075 ( .A(n1014), .B(n1015), .C(n1016), .Y(n773) );
  OR2XL U1076 ( .A(n559), .B(n560), .Y(n537) );
  NAND2X2 U1077 ( .A(n985), .B(n523), .Y(n455) );
  INVX1 U1078 ( .A(n996), .Y(n1098) );
  CLKBUFX3 U1079 ( .A(n409), .Y(n1039) );
  OAI32XL U1080 ( .A0(n456), .A1(n1102), .A2(n1101), .B0(n1108), .B1(n1106), 
        .Y(n409) );
  CLKINVX1 U1081 ( .A(n413), .Y(n1100) );
  NOR2X2 U1082 ( .A(n547), .B(n1085), .Y(n528) );
  NAND2X1 U1083 ( .A(n541), .B(n531), .Y(n532) );
  CLKINVX1 U1084 ( .A(n547), .Y(n1086) );
  NAND2X1 U1085 ( .A(n1105), .B(n980), .Y(n559) );
  NAND2X1 U1086 ( .A(n1096), .B(n489), .Y(n545) );
  NAND2XL U1087 ( .A(n996), .B(n339), .Y(n560) );
  NAND2X1 U1088 ( .A(n328), .B(n1050), .Y(n329) );
  CLKBUFX3 U1089 ( .A(n316), .Y(n1056) );
  CLKBUFX3 U1090 ( .A(n316), .Y(n1055) );
  CLKBUFX3 U1091 ( .A(n314), .Y(n1059) );
  CLKBUFX3 U1092 ( .A(n313), .Y(n1061) );
  CLKBUFX3 U1093 ( .A(n318), .Y(n1051) );
  CLKBUFX3 U1095 ( .A(n315), .Y(n1057) );
  CLKBUFX3 U1096 ( .A(n1045), .Y(n1046) );
  CLKBUFX3 U1097 ( .A(n1045), .Y(n1048) );
  CLKBUFX3 U1098 ( .A(n1045), .Y(n1047) );
  OAI222XL U1099 ( .A0(n1160), .A1(n422), .B0(n486), .B1(n916), .C0(n1153), 
        .C1(n1037), .Y(n841) );
  OAI222XL U1100 ( .A0(n1141), .A1(n422), .B0(n396), .B1(n916), .C0(n1134), 
        .C1(n1037), .Y(n774) );
  OAI222XL U1101 ( .A0(n1120), .A1(n422), .B0(n398), .B1(n916), .C0(n1121), 
        .C1(n1037), .Y(n775) );
  CLKINVX1 U1102 ( .A(n526), .Y(n1097) );
  CLKINVX1 U1103 ( .A(n459), .Y(n1101) );
  CLKINVX1 U1104 ( .A(n383), .Y(n1109) );
  OAI211X1 U1105 ( .A0(n1044), .A1(n487), .B0(n488), .C0(n422), .Y(n424) );
  OR2X1 U1106 ( .A(n460), .B(n1097), .Y(n515) );
  CLKBUFX3 U1107 ( .A(n403), .Y(n1041) );
  OAI32XL U1108 ( .A0(n456), .A1(n1101), .A2(n457), .B0(n458), .B1(n1106), .Y(
        n403) );
  CLKBUFX3 U1109 ( .A(n428), .Y(n1034) );
  NOR3X1 U1110 ( .A(n513), .B(n1093), .C(n512), .Y(n428) );
  NAND2X1 U1111 ( .A(n562), .B(n384), .Y(n339) );
  CLKINVX1 U1112 ( .A(n512), .Y(n1094) );
  NAND3X1 U1113 ( .A(n1087), .B(n488), .C(n522), .Y(n549) );
  OAI21XL U1114 ( .A0(n543), .A1(n1087), .B0(n489), .Y(n542) );
  CLKINVX1 U1115 ( .A(n421), .Y(n1110) );
  OAI22XL U1116 ( .A0(n1092), .A1(n486), .B0(n1160), .B1(n1033), .Y(n842) );
  OAI22XL U1117 ( .A0(n1213), .A1(n1033), .B0(n1092), .B1(n439), .Y(n780) );
  OAI22XL U1118 ( .A0(n1205), .A1(n1033), .B0(n1092), .B1(n441), .Y(n782) );
  OAI22XL U1119 ( .A0(n1198), .A1(n1033), .B0(n1092), .B1(n443), .Y(n784) );
  OAI22XL U1120 ( .A0(n956), .A1(n1033), .B0(n1092), .B1(n445), .Y(n786) );
  OAI22XL U1121 ( .A0(n1183), .A1(n1033), .B0(n1092), .B1(n447), .Y(n788) );
  OAI22XL U1122 ( .A0(n1175), .A1(n1033), .B0(n1092), .B1(n449), .Y(n790) );
  OAI22XL U1123 ( .A0(n1167), .A1(n1033), .B0(n1092), .B1(n451), .Y(n792) );
  OAI22XL U1124 ( .A0(n1149), .A1(n1033), .B0(n1092), .B1(n400), .Y(n751) );
  OAI22XL U1125 ( .A0(n1141), .A1(n1033), .B0(n1092), .B1(n396), .Y(n747) );
  OAI22XL U1126 ( .A0(n1133), .A1(n1033), .B0(n1092), .B1(n392), .Y(n745) );
  OAI22XL U1127 ( .A0(n1120), .A1(n1033), .B0(n1092), .B1(n398), .Y(n749) );
  CLKINVX1 U1128 ( .A(n461), .Y(n1099) );
  CLKBUFX3 U1129 ( .A(n406), .Y(n1040) );
  OAI32XL U1130 ( .A0(n456), .A1(n1102), .A2(n459), .B0(n460), .B1(n1106), .Y(
        n406) );
  NOR3X1 U1131 ( .A(n512), .B(n513), .C(n514), .Y(n429) );
  CLKBUFX3 U1132 ( .A(n319), .Y(n1043) );
  OAI31XL U1133 ( .A0(n322), .A1(n1050), .A2(n323), .B0(n324), .Y(n319) );
  OR3X2 U1134 ( .A(n325), .B(n326), .C(n327), .Y(n322) );
  AND2X2 U1135 ( .A(n324), .B(n488), .Y(n541) );
  NOR2BX2 U1136 ( .AN(n382), .B(n381), .Y(n352) );
  NOR2BX2 U1137 ( .AN(n381), .B(n382), .Y(n351) );
  OAI21X1 U1138 ( .A0(n332), .A1(n1002), .B0(n1050), .Y(n328) );
  AOI32X1 U1139 ( .A0(n572), .A1(n1087), .A2(n1097), .B0(n564), .B1(n526), .Y(
        n570) );
  NAND2X2 U1140 ( .A(n381), .B(n382), .Y(n347) );
  NOR2X1 U1141 ( .A(n522), .B(n566), .Y(n567) );
  NAND2X1 U1142 ( .A(n546), .B(n526), .Y(n489) );
  CLKINVX1 U1143 ( .A(n539), .Y(n1105) );
  OA21XL U1144 ( .A0(n518), .A1(n980), .B0(n1105), .Y(n556) );
  CLKINVX1 U1145 ( .A(n521), .Y(n1096) );
  CLKINVX1 U1146 ( .A(n332), .Y(n1111) );
  CLKBUFX3 U1147 ( .A(n1084), .Y(n1045) );
  CLKINVX1 U1148 ( .A(N386), .Y(n1083) );
  CLKINVX1 U1149 ( .A(N378), .Y(n1072) );
  MXI2X2 U1150 ( .A(n106), .B(n1074), .S0(net5660), .Y(n888) );
  CLKINVX1 U1151 ( .A(N394), .Y(n1074) );
  CLKMX2X4 U1152 ( .A(CNT3[1]), .B(N395), .S0(net5660), .Y(n887) );
  CLKMX2X4 U1153 ( .A(CNT3[2]), .B(N396), .S0(net5660), .Y(n886) );
  CLKMX2X4 U1154 ( .A(CNT3[3]), .B(N397), .S0(net5660), .Y(n885) );
  CLKMX2X4 U1155 ( .A(CNT3[4]), .B(N398), .S0(net5660), .Y(n884) );
  CLKMX2X4 U1156 ( .A(CNT3[5]), .B(N399), .S0(net5660), .Y(n883) );
  CLKMX2X4 U1157 ( .A(CNT3[6]), .B(N400), .S0(net5660), .Y(n882) );
  INVX1 U1158 ( .A(N402), .Y(n1075) );
  CLKINVX1 U1159 ( .A(N418), .Y(n1073) );
  AOI211X1 U1160 ( .A0(cs[0]), .A1(n575), .B0(n576), .C0(n567), .Y(n574) );
  NAND2X1 U1161 ( .A(n555), .B(n1105), .Y(n576) );
  OAI2BB1X1 U1162 ( .A0N(n573), .A1N(n384), .B0(n570), .Y(n575) );
  NOR2BX1 U1163 ( .AN(n568), .B(n569), .Y(n863) );
  OAI222X4 U1164 ( .A0(n260), .A1(n517), .B0(n252), .B1(n515), .C0(n520), .C1(
        n487), .Y(n514) );
  XNOR2X1 U1165 ( .A(N488), .B(n1044), .Y(n520) );
  CLKINVX1 U1166 ( .A(\ListB[1][5] ), .Y(n1200) );
  CLKINVX1 U1168 ( .A(\ListB[1][4] ), .Y(n1193) );
  CLKINVX1 U1170 ( .A(\ListB[1][3] ), .Y(n1186) );
  CLKINVX1 U1172 ( .A(\ListB[1][2] ), .Y(n1178) );
  CLKINVX1 U1174 ( .A(\ListB[1][1] ), .Y(n1170) );
  CLKINVX1 U1176 ( .A(\ListB[1][0] ), .Y(n1162) );
  CLKINVX1 U1180 ( .A(\ListB[5][6] ), .Y(n1212) );
  CLKINVX1 U1181 ( .A(\ListB[5][7] ), .Y(n1158) );
  CLKINVX1 U1182 ( .A(\ListB[1][6] ), .Y(n1208) );
  CLKINVX1 U1183 ( .A(\ListB[1][7] ), .Y(n1154) );
  OAI222XL U1184 ( .A0(n440), .A1(n982), .B0(n918), .B1(n92), .C0(n1031), .C1(
        n1211), .Y(n819) );
  CLKINVX1 U1185 ( .A(\ListB[4][6] ), .Y(n1211) );
  OAI222XL U1186 ( .A0(n440), .A1(n981), .B0(n993), .B1(n84), .C0(n1039), .C1(
        n1210), .Y(n811) );
  CLKINVX1 U1187 ( .A(\ListB[3][6] ), .Y(n1210) );
  OAI222XL U1188 ( .A0(n442), .A1(n982), .B0(n918), .B1(n93), .C0(n1031), .C1(
        n1203), .Y(n820) );
  CLKINVX1 U1189 ( .A(\ListB[4][5] ), .Y(n1203) );
  OAI222XL U1190 ( .A0(n442), .A1(n981), .B0(n993), .B1(n85), .C0(n1039), .C1(
        n1202), .Y(n812) );
  CLKINVX1 U1191 ( .A(\ListB[3][5] ), .Y(n1202) );
  OAI222XL U1192 ( .A0(n444), .A1(n982), .B0(n918), .B1(n94), .C0(n1031), .C1(
        n1196), .Y(n821) );
  CLKINVX1 U1193 ( .A(\ListB[4][4] ), .Y(n1196) );
  OAI222XL U1194 ( .A0(n444), .A1(n981), .B0(n993), .B1(n86), .C0(n1039), .C1(
        n1195), .Y(n813) );
  CLKINVX1 U1195 ( .A(\ListB[3][4] ), .Y(n1195) );
  OAI222XL U1196 ( .A0(n446), .A1(n982), .B0(n918), .B1(n95), .C0(n1031), .C1(
        n1189), .Y(n822) );
  CLKINVX1 U1197 ( .A(\ListB[4][3] ), .Y(n1189) );
  OAI222XL U1198 ( .A0(n446), .A1(n981), .B0(n993), .B1(n87), .C0(n1039), .C1(
        n1188), .Y(n814) );
  CLKINVX1 U1199 ( .A(\ListB[3][3] ), .Y(n1188) );
  OAI222XL U1200 ( .A0(n448), .A1(n982), .B0(n918), .B1(n96), .C0(n1031), .C1(
        n1181), .Y(n823) );
  CLKINVX1 U1201 ( .A(\ListB[4][2] ), .Y(n1181) );
  OAI222XL U1202 ( .A0(n448), .A1(n981), .B0(n993), .B1(n88), .C0(n1039), .C1(
        n1180), .Y(n815) );
  CLKINVX1 U1203 ( .A(\ListB[3][2] ), .Y(n1180) );
  OAI222XL U1204 ( .A0(n450), .A1(n982), .B0(n918), .B1(n97), .C0(n1031), .C1(
        n1173), .Y(n824) );
  CLKINVX1 U1205 ( .A(\ListB[4][1] ), .Y(n1173) );
  OAI222XL U1206 ( .A0(n450), .A1(n981), .B0(n993), .B1(n89), .C0(n1039), .C1(
        n1172), .Y(n816) );
  CLKINVX1 U1207 ( .A(\ListB[3][1] ), .Y(n1172) );
  OAI222XL U1208 ( .A0(n452), .A1(n982), .B0(n918), .B1(n98), .C0(n1031), .C1(
        n1165), .Y(n825) );
  CLKINVX1 U1209 ( .A(\ListB[4][0] ), .Y(n1165) );
  OAI222XL U1210 ( .A0(n452), .A1(n981), .B0(n993), .B1(n90), .C0(n1039), .C1(
        n1164), .Y(n817) );
  CLKINVX1 U1211 ( .A(\ListB[3][0] ), .Y(n1164) );
  CLKINVX1 U1212 ( .A(\ListB[4][7] ), .Y(n1157) );
  CLKINVX1 U1213 ( .A(\ListB[3][7] ), .Y(n1156) );
  AND2X2 U1214 ( .A(n472), .B(n473), .Y(n439) );
  AOI222XL U1215 ( .A0(\ListB[2][6] ), .A1(n1000), .B0(\ListB[4][6] ), .B1(
        n1001), .C0(\ListB[3][6] ), .C1(n988), .Y(n472) );
  AOI222XL U1216 ( .A0(\ListB[5][6] ), .A1(n987), .B0(\ListB[1][6] ), .B1(
        n1034), .C0(\ListB[0][6] ), .C1(n1035), .Y(n473) );
  AND2X2 U1217 ( .A(n474), .B(n475), .Y(n441) );
  AOI222XL U1218 ( .A0(\ListB[2][5] ), .A1(n1000), .B0(\ListB[4][5] ), .B1(
        n1001), .C0(\ListB[3][5] ), .C1(n988), .Y(n474) );
  AOI222XL U1219 ( .A0(\ListB[5][5] ), .A1(n987), .B0(\ListB[1][5] ), .B1(
        n1034), .C0(\ListB[0][5] ), .C1(n1035), .Y(n475) );
  AND2X2 U1220 ( .A(n476), .B(n477), .Y(n443) );
  AOI222XL U1221 ( .A0(\ListB[2][4] ), .A1(n1000), .B0(\ListB[4][4] ), .B1(
        n1001), .C0(\ListB[3][4] ), .C1(n988), .Y(n476) );
  AOI222XL U1222 ( .A0(\ListB[5][4] ), .A1(n987), .B0(\ListB[1][4] ), .B1(
        n1034), .C0(\ListB[0][4] ), .C1(n1035), .Y(n477) );
  AND2X2 U1223 ( .A(n478), .B(n479), .Y(n445) );
  AOI222XL U1224 ( .A0(\ListB[2][3] ), .A1(n1000), .B0(\ListB[4][3] ), .B1(
        n1001), .C0(\ListB[3][3] ), .C1(n988), .Y(n478) );
  AOI222XL U1225 ( .A0(\ListB[5][3] ), .A1(n987), .B0(\ListB[1][3] ), .B1(
        n1034), .C0(\ListB[0][3] ), .C1(n1035), .Y(n479) );
  AND2X2 U1226 ( .A(n480), .B(n481), .Y(n447) );
  AOI222XL U1227 ( .A0(\ListB[2][2] ), .A1(n1000), .B0(\ListB[4][2] ), .B1(
        n1001), .C0(\ListB[3][2] ), .C1(n988), .Y(n480) );
  AOI222XL U1228 ( .A0(\ListB[5][2] ), .A1(n987), .B0(\ListB[1][2] ), .B1(
        n1034), .C0(\ListB[0][2] ), .C1(n1035), .Y(n481) );
  AND2X2 U1229 ( .A(n482), .B(n483), .Y(n449) );
  AOI222XL U1230 ( .A0(\ListB[2][1] ), .A1(n1000), .B0(\ListB[4][1] ), .B1(
        n1001), .C0(\ListB[3][1] ), .C1(n988), .Y(n482) );
  AOI222XL U1231 ( .A0(\ListB[5][1] ), .A1(n987), .B0(\ListB[1][1] ), .B1(
        n1034), .C0(\ListB[0][1] ), .C1(n1035), .Y(n483) );
  AOI222XL U1232 ( .A0(\ListB[2][0] ), .A1(n1000), .B0(\ListB[4][0] ), .B1(
        n1001), .C0(\ListB[3][0] ), .C1(n988), .Y(n484) );
  AOI222XL U1233 ( .A0(\ListB[5][0] ), .A1(n987), .B0(\ListB[1][0] ), .B1(
        n1034), .C0(\ListB[0][0] ), .C1(n1035), .Y(n485) );
  AND2X2 U1234 ( .A(n510), .B(n511), .Y(n486) );
  AOI222XL U1235 ( .A0(\ListB[2][7] ), .A1(n1000), .B0(\ListB[4][7] ), .B1(
        n1001), .C0(\ListB[3][7] ), .C1(n988), .Y(n510) );
  AOI222XL U1236 ( .A0(\ListB[5][7] ), .A1(n987), .B0(\ListB[1][7] ), .B1(
        n1034), .C0(\ListB[0][7] ), .C1(n1035), .Y(n511) );
  AOI222XL U1237 ( .A0(\ListA[2][0] ), .A1(n1000), .B0(\ListA[4][0] ), .B1(
        n1001), .C0(\ListA[3][0] ), .C1(n988), .Y(n437) );
  AOI222XL U1238 ( .A0(\ListA[5][0] ), .A1(n987), .B0(\ListA[1][0] ), .B1(
        n1034), .C0(\ListA[0][0] ), .C1(n1035), .Y(n438) );
  AND2X2 U1239 ( .A(n433), .B(n434), .Y(n396) );
  AOI222XL U1240 ( .A0(\ListA[2][2] ), .A1(n1000), .B0(\ListA[4][2] ), .B1(
        n1001), .C0(\ListA[3][2] ), .C1(n988), .Y(n433) );
  AOI222XL U1241 ( .A0(\ListA[5][2] ), .A1(n987), .B0(\ListA[1][2] ), .B1(
        n1034), .C0(\ListA[0][2] ), .C1(n1035), .Y(n434) );
  AOI222XL U1242 ( .A0(\ListA[2][3] ), .A1(n1000), .B0(\ListA[4][3] ), .B1(
        n1001), .C0(\ListA[3][3] ), .C1(n988), .Y(n425) );
  AOI222XL U1243 ( .A0(\ListA[5][3] ), .A1(n987), .B0(\ListA[1][3] ), .B1(
        n1034), .C0(\ListA[0][3] ), .C1(n1035), .Y(n426) );
  AND2X2 U1244 ( .A(n435), .B(n436), .Y(n398) );
  AOI222XL U1245 ( .A0(\ListA[2][1] ), .A1(n1000), .B0(\ListA[4][1] ), .B1(
        n1001), .C0(\ListA[3][1] ), .C1(n988), .Y(n435) );
  AOI222XL U1246 ( .A0(\ListA[5][1] ), .A1(n987), .B0(\ListA[1][1] ), .B1(
        n1034), .C0(\ListA[0][1] ), .C1(n1035), .Y(n436) );
  OAI221XL U1247 ( .A0(n401), .A1(n982), .B0(n1147), .B1(n1031), .C0(n918), 
        .Y(n768) );
  CLKINVX1 U1248 ( .A(\ListA[4][0] ), .Y(n1147) );
  OAI221XL U1249 ( .A0(n397), .A1(n982), .B0(n1139), .B1(n1031), .C0(n918), 
        .Y(n766) );
  CLKINVX1 U1250 ( .A(\ListA[4][2] ), .Y(n1139) );
  OAI2BB2XL U1251 ( .B0(n394), .B1(n982), .A0N(\ListA[4][3] ), .A1N(n413), .Y(
        n765) );
  NOR3X1 U1252 ( .A(n458), .B(cnt2[1]), .C(n1097), .Y(n521) );
  OAI22XL U1253 ( .A0(n246), .A1(n1037), .B0(n258), .B1(n422), .Y(n777) );
  OAI2BB2XL U1254 ( .B0(n399), .B1(n982), .A0N(\ListA[4][1] ), .A1N(n413), .Y(
        n767) );
  OAI22XL U1255 ( .A0(n247), .A1(n1037), .B0(n259), .B1(n422), .Y(n778) );
  OAI22XL U1256 ( .A0(n248), .A1(n1037), .B0(n260), .B1(n422), .Y(n779) );
  CLKBUFX3 U1257 ( .A(n415), .Y(n1038) );
  OAI31XL U1258 ( .A0(n457), .A1(n1101), .A2(n1099), .B0(n470), .Y(n415) );
  NAND4XL U1259 ( .A(n1010), .B(cnt[2]), .C(n1044), .D(n140), .Y(n470) );
  AOI221X4 U1260 ( .A0(n985), .A1(RegA_t[3]), .B0(RegB_t[3]), .B1(n1098), .C0(
        n418), .Y(n394) );
  OA21XL U1261 ( .A0(n1110), .A1(n253), .B0(n999), .Y(n418) );
  AOI222X4 U1262 ( .A0(n421), .A1(n999), .B0(n985), .B1(RegA_t[1]), .C0(
        RegB_t[1]), .C1(n1098), .Y(n399) );
  AOI222X4 U1263 ( .A0(N488), .A1(n999), .B0(n985), .B1(RegA_t[0]), .C0(
        RegB_t[0]), .C1(n1098), .Y(n401) );
  AOI221X4 U1264 ( .A0(n985), .A1(RegA_t[2]), .B0(RegB_t[2]), .B1(n1098), .C0(
        n420), .Y(n397) );
  AOI2BB2X1 U1265 ( .B0(n1036), .B1(RegB_t[0]), .A0N(n1036), .A1N(n1142), .Y(
        n385) );
  AOI2BB2X1 U1266 ( .B0(n1036), .B1(RegA_t[0]), .A0N(n1149), .A1N(n1036), .Y(
        n369) );
  AOI2BB2X1 U1267 ( .B0(n1036), .B1(RegB_t[2]), .A0N(n1134), .A1N(n1036), .Y(
        n375) );
  AOI2BB2X1 U1268 ( .B0(n1036), .B1(RegA_t[2]), .A0N(n1141), .A1N(n1036), .Y(
        n363) );
  AOI2BB2X1 U1269 ( .B0(n1036), .B1(RegB_t[3]), .A0N(n1127), .A1N(n1036), .Y(
        n372) );
  AOI2BB2X1 U1270 ( .B0(n1036), .B1(RegA_t[3]), .A0N(n1133), .A1N(n1036), .Y(
        n354) );
  AOI2BB2X1 U1271 ( .B0(n1036), .B1(RegB_t[1]), .A0N(n1121), .A1N(n1036), .Y(
        n378) );
  AOI2BB2X1 U1272 ( .B0(n1036), .B1(RegA_t[1]), .A0N(n1120), .A1N(n1036), .Y(
        n366) );
  OAI211X1 U1273 ( .A0(n340), .A1(n341), .B0(n149), .C0(n342), .Y(n321) );
  NOR4X1 U1274 ( .A(n343), .B(n344), .C(n345), .D(n346), .Y(n340) );
  NOR4X1 U1275 ( .A(n326), .B(n325), .C(n327), .D(n323), .Y(n341) );
  OAI222XL U1276 ( .A0(n440), .A1(n983), .B0(n992), .B1(n100), .C0(n1040), 
        .C1(n1209), .Y(n803) );
  CLKINVX1 U1277 ( .A(\ListB[2][6] ), .Y(n1209) );
  OAI222XL U1278 ( .A0(n442), .A1(n997), .B0(n998), .B1(n109), .C0(n1038), 
        .C1(n1204), .Y(n828) );
  CLKINVX1 U1279 ( .A(\ListB[5][5] ), .Y(n1204) );
  OAI222XL U1280 ( .A0(n442), .A1(n983), .B0(n992), .B1(n101), .C0(n1040), 
        .C1(n1201), .Y(n804) );
  CLKINVX1 U1281 ( .A(\ListB[2][5] ), .Y(n1201) );
  OAI222XL U1282 ( .A0(n444), .A1(n997), .B0(n998), .B1(n110), .C0(n1038), 
        .C1(n1197), .Y(n829) );
  CLKINVX1 U1283 ( .A(\ListB[5][4] ), .Y(n1197) );
  OAI222XL U1284 ( .A0(n444), .A1(n983), .B0(n992), .B1(n102), .C0(n1040), 
        .C1(n1194), .Y(n805) );
  CLKINVX1 U1285 ( .A(\ListB[2][4] ), .Y(n1194) );
  OAI222XL U1286 ( .A0(n446), .A1(n997), .B0(n998), .B1(n111), .C0(n1038), 
        .C1(n1190), .Y(n830) );
  CLKINVX1 U1287 ( .A(\ListB[5][3] ), .Y(n1190) );
  OAI222XL U1288 ( .A0(n446), .A1(n983), .B0(n992), .B1(n103), .C0(n1040), 
        .C1(n1187), .Y(n806) );
  CLKINVX1 U1289 ( .A(\ListB[2][3] ), .Y(n1187) );
  OAI222XL U1290 ( .A0(n448), .A1(n997), .B0(n998), .B1(n112), .C0(n1038), 
        .C1(n1182), .Y(n831) );
  CLKINVX1 U1291 ( .A(\ListB[5][2] ), .Y(n1182) );
  OAI222XL U1292 ( .A0(n448), .A1(n983), .B0(n992), .B1(n104), .C0(n1040), 
        .C1(n1179), .Y(n807) );
  CLKINVX1 U1293 ( .A(\ListB[2][2] ), .Y(n1179) );
  OAI222XL U1294 ( .A0(n450), .A1(n997), .B0(n998), .B1(n113), .C0(n1038), 
        .C1(n1174), .Y(n832) );
  CLKINVX1 U1295 ( .A(\ListB[5][1] ), .Y(n1174) );
  OAI222XL U1296 ( .A0(n450), .A1(n983), .B0(n992), .B1(n105), .C0(n1040), 
        .C1(n1171), .Y(n808) );
  CLKINVX1 U1297 ( .A(\ListB[2][1] ), .Y(n1171) );
  OAI222XL U1298 ( .A0(n452), .A1(n997), .B0(n998), .B1(n114), .C0(n1038), 
        .C1(n1166), .Y(n833) );
  CLKINVX1 U1299 ( .A(\ListB[5][0] ), .Y(n1166) );
  OAI222XL U1300 ( .A0(n452), .A1(n983), .B0(n992), .B1(n106), .C0(n1040), 
        .C1(n1163), .Y(n809) );
  CLKINVX1 U1301 ( .A(\ListB[2][0] ), .Y(n1163) );
  CLKINVX1 U1302 ( .A(\ListB[2][7] ), .Y(n1155) );
  OAI32X1 U1303 ( .A0(n530), .A1(int_i[2]), .A2(n259), .B0(n540), .B1(n258), 
        .Y(n851) );
  OA21XL U1304 ( .A0(int_i[1]), .A1(n531), .B0(n529), .Y(n540) );
  OAI221XL U1305 ( .A0(n399), .A1(n983), .B0(n1125), .B1(n1040), .C0(n992), 
        .Y(n759) );
  CLKINVX1 U1306 ( .A(\ListA[2][1] ), .Y(n1125) );
  OAI221XL U1307 ( .A0(n399), .A1(n997), .B0(n1124), .B1(n1038), .C0(n998), 
        .Y(n771) );
  CLKINVX1 U1308 ( .A(\ListA[5][1] ), .Y(n1124) );
  OAI221XL U1309 ( .A0(n399), .A1(n984), .B0(n1122), .B1(n1041), .C0(n994), 
        .Y(n755) );
  CLKINVX1 U1310 ( .A(\ListA[1][1] ), .Y(n1122) );
  OAI221XL U1311 ( .A0(n401), .A1(n983), .B0(n1145), .B1(n1040), .C0(n992), 
        .Y(n760) );
  CLKINVX1 U1312 ( .A(\ListA[2][0] ), .Y(n1145) );
  OAI221XL U1313 ( .A0(n401), .A1(n991), .B0(n1032), .B1(n1143), .C0(n995), 
        .Y(n752) );
  CLKINVX1 U1314 ( .A(\ListA[0][0] ), .Y(n1143) );
  XOR2X1 U1315 ( .A(n253), .B(n563), .Y(n518) );
  OAI221XL U1316 ( .A0(n397), .A1(n997), .B0(n1140), .B1(n1038), .C0(n998), 
        .Y(n770) );
  CLKINVX1 U1317 ( .A(\ListA[5][2] ), .Y(n1140) );
  OAI221XL U1318 ( .A0(n397), .A1(n981), .B0(n1138), .B1(n1039), .C0(n993), 
        .Y(n762) );
  CLKINVX1 U1319 ( .A(\ListA[3][2] ), .Y(n1138) );
  OAI22XL U1320 ( .A0(n1132), .A1(n1038), .B0(n394), .B1(n997), .Y(n769) );
  CLKINVX1 U1321 ( .A(\ListA[5][3] ), .Y(n1132) );
  OAI22XL U1322 ( .A0(n1131), .A1(n1039), .B0(n394), .B1(n981), .Y(n761) );
  CLKINVX1 U1323 ( .A(\ListA[3][3] ), .Y(n1131) );
  OAI22XL U1324 ( .A0(n1130), .A1(n1040), .B0(n394), .B1(n983), .Y(n757) );
  CLKINVX1 U1325 ( .A(\ListA[2][3] ), .Y(n1130) );
  OAI22XL U1326 ( .A0(n1129), .A1(n1041), .B0(n394), .B1(n984), .Y(n753) );
  CLKINVX1 U1327 ( .A(\ListA[1][3] ), .Y(n1129) );
  OAI22XL U1328 ( .A0(n1128), .A1(n1032), .B0(n394), .B1(n991), .Y(n746) );
  CLKINVX1 U1329 ( .A(\ListA[0][3] ), .Y(n1128) );
  OAI22XL U1330 ( .A0(n1032), .A1(n1126), .B0(n399), .B1(n991), .Y(n750) );
  CLKINVX1 U1331 ( .A(\ListA[0][1] ), .Y(n1126) );
  OAI22XL U1332 ( .A0(n1123), .A1(n1039), .B0(n399), .B1(n981), .Y(n763) );
  CLKINVX1 U1333 ( .A(\ListA[3][1] ), .Y(n1123) );
  OAI22XL U1334 ( .A0(n1148), .A1(n1038), .B0(n401), .B1(n997), .Y(n772) );
  CLKINVX1 U1335 ( .A(\ListA[5][0] ), .Y(n1148) );
  OAI22XL U1336 ( .A0(n1146), .A1(n1039), .B0(n401), .B1(n981), .Y(n764) );
  CLKINVX1 U1337 ( .A(\ListA[3][0] ), .Y(n1146) );
  OAI22XL U1338 ( .A0(n1144), .A1(n1041), .B0(n401), .B1(n984), .Y(n756) );
  CLKINVX1 U1339 ( .A(\ListA[1][0] ), .Y(n1144) );
  OAI22XL U1340 ( .A0(n1137), .A1(n1040), .B0(n397), .B1(n983), .Y(n758) );
  CLKINVX1 U1341 ( .A(\ListA[2][2] ), .Y(n1137) );
  OAI22XL U1342 ( .A0(n1136), .A1(n1041), .B0(n397), .B1(n984), .Y(n754) );
  CLKINVX1 U1343 ( .A(\ListA[1][2] ), .Y(n1136) );
  OAI22XL U1344 ( .A0(n1032), .A1(n1135), .B0(n397), .B1(n991), .Y(n748) );
  CLKINVX1 U1345 ( .A(\ListA[0][2] ), .Y(n1135) );
  NOR2X1 U1346 ( .A(n543), .B(cnt[2]), .Y(n525) );
  OAI2BB2XL U1347 ( .B0(n282), .B1(n1043), .A0N(N718), .A1N(n320), .Y(n595) );
  OAI2BB2XL U1348 ( .B0(n363), .B1(n1006), .A0N(n1006), .A1N(\Tree_0[1][2] ), 
        .Y(n720) );
  OAI2BB2XL U1349 ( .B0(n363), .B1(n1007), .A0N(n1007), .A1N(\Tree_0[2][2] ), 
        .Y(n719) );
  OAI2BB2XL U1350 ( .B0(n363), .B1(n1042), .A0N(n1042), .A1N(\Tree_0[4][2] ), 
        .Y(n718) );
  OAI2BB2XL U1351 ( .B0(n369), .B1(n1006), .A0N(n1006), .A1N(\Tree_0[1][0] ), 
        .Y(n728) );
  OAI2BB2XL U1352 ( .B0(n369), .B1(n1007), .A0N(n1007), .A1N(\Tree_0[2][0] ), 
        .Y(n727) );
  OAI2BB2XL U1353 ( .B0(n369), .B1(n1042), .A0N(n1042), .A1N(\Tree_0[4][0] ), 
        .Y(n726) );
  OAI2BB2XL U1354 ( .B0(n375), .B1(n1006), .A0N(n1006), .A1N(\Tree_1[1][2] ), 
        .Y(n736) );
  OAI2BB2XL U1355 ( .B0(n375), .B1(n1007), .A0N(n1007), .A1N(\Tree_1[2][2] ), 
        .Y(n735) );
  OAI2BB2XL U1356 ( .B0(n375), .B1(n1042), .A0N(n1042), .A1N(\Tree_1[4][2] ), 
        .Y(n734) );
  OAI2BB2XL U1357 ( .B0(n378), .B1(n1006), .A0N(n1006), .A1N(\Tree_1[1][1] ), 
        .Y(n740) );
  OAI2BB2XL U1358 ( .B0(n378), .B1(n1007), .A0N(n1007), .A1N(\Tree_1[2][1] ), 
        .Y(n739) );
  OAI2BB2XL U1359 ( .B0(n378), .B1(n1042), .A0N(n1042), .A1N(\Tree_1[4][1] ), 
        .Y(n738) );
  OAI2BB2XL U1360 ( .B0(n366), .B1(n1006), .A0N(n1006), .A1N(\Tree_0[1][1] ), 
        .Y(n724) );
  OAI2BB2XL U1361 ( .B0(n366), .B1(n1007), .A0N(n1007), .A1N(\Tree_0[2][1] ), 
        .Y(n723) );
  OAI2BB2XL U1362 ( .B0(n366), .B1(n1042), .A0N(n1042), .A1N(\Tree_0[4][1] ), 
        .Y(n722) );
  OAI2BB2XL U1363 ( .B0(n372), .B1(n1006), .A0N(n1006), .A1N(\Tree_1[1][3] ), 
        .Y(n732) );
  OAI2BB2XL U1364 ( .B0(n372), .B1(n1007), .A0N(n1007), .A1N(\Tree_1[2][3] ), 
        .Y(n731) );
  OAI2BB2XL U1365 ( .B0(n372), .B1(n1042), .A0N(n1042), .A1N(\Tree_1[4][3] ), 
        .Y(n730) );
  OAI2BB2XL U1366 ( .B0(n354), .B1(n1006), .A0N(n1006), .A1N(\Tree_0[1][3] ), 
        .Y(n716) );
  OAI2BB2XL U1367 ( .B0(n354), .B1(n1007), .A0N(n1007), .A1N(\Tree_0[2][3] ), 
        .Y(n715) );
  OAI2BB2XL U1368 ( .B0(n354), .B1(n1042), .A0N(n1042), .A1N(\Tree_0[4][3] ), 
        .Y(n714) );
  OAI2BB2XL U1369 ( .B0(n385), .B1(n1006), .A0N(n1006), .A1N(\Tree_1[1][0] ), 
        .Y(n744) );
  OAI2BB2XL U1370 ( .B0(n385), .B1(n1007), .A0N(n1007), .A1N(\Tree_1[2][0] ), 
        .Y(n743) );
  OAI2BB2XL U1371 ( .B0(n385), .B1(n1042), .A0N(n1042), .A1N(\Tree_1[4][0] ), 
        .Y(n742) );
  OAI2BB2XL U1372 ( .B0(n1043), .B1(n281), .A0N(N719), .A1N(n320), .Y(n644) );
  OAI2BB2XL U1373 ( .B0(n1043), .B1(n283), .A0N(N717), .A1N(n320), .Y(n602) );
  OAI2BB2XL U1374 ( .B0(n1043), .B1(n284), .A0N(N716), .A1N(n320), .Y(n609) );
  OAI2BB2XL U1375 ( .B0(n1043), .B1(n285), .A0N(N715), .A1N(n320), .Y(n616) );
  OAI2BB2XL U1376 ( .B0(n1043), .B1(n286), .A0N(N714), .A1N(n320), .Y(n623) );
  OAI2BB2XL U1377 ( .B0(n1043), .B1(n287), .A0N(N713), .A1N(n320), .Y(n630) );
  OAI2BB2XL U1378 ( .B0(n1043), .B1(n288), .A0N(N712), .A1N(n320), .Y(n637) );
  OR2X1 U1379 ( .A(n522), .B(cnt[1]), .Y(n487) );
  OA21XL U1380 ( .A0(int_i[0]), .A1(n531), .B0(n532), .Y(n529) );
  NOR2X1 U1381 ( .A(n140), .B(n1087), .Y(n342) );
  AO22X1 U1382 ( .A0(cnt[6]), .A1(n528), .B0(N446), .B1(n1085), .Y(n857) );
  AO22X1 U1383 ( .A0(cnt[5]), .A1(n528), .B0(N445), .B1(n1085), .Y(n844) );
  AO22X1 U1384 ( .A0(cnt[4]), .A1(n528), .B0(N444), .B1(n1085), .Y(n845) );
  AO22X1 U1385 ( .A0(cnt[3]), .A1(n528), .B0(N443), .B1(n1085), .Y(n846) );
  NOR4X1 U1386 ( .A(cnt[3]), .B(cnt[4]), .C(cnt[5]), .D(cnt[6]), .Y(n577) );
  OAI222XL U1387 ( .A0(int_i[0]), .A1(n1050), .B0(n252), .B1(n329), .C0(n1152), 
        .C1(n328), .Y(n648) );
  OAI222XL U1388 ( .A0(n251), .A1(n329), .B0(n333), .B1(n1050), .C0(n1151), 
        .C1(n328), .Y(n647) );
  OAI222XL U1389 ( .A0(n249), .A1(n329), .B0(n330), .B1(n1050), .C0(n1150), 
        .C1(n328), .Y(n646) );
  XNOR2X1 U1390 ( .A(n277), .B(tmp_T1[3]), .Y(n323) );
  XOR2X1 U1391 ( .A(node[2]), .B(tmp_T1[2]), .Y(n327) );
  XOR2X1 U1392 ( .A(node[0]), .B(tmp_T1[0]), .Y(n326) );
  XOR2X1 U1393 ( .A(node[1]), .B(tmp_T1[1]), .Y(n325) );
  OAI221XL U1394 ( .A0(int_j[1]), .A1(n533), .B0(n534), .B1(n251), .C0(n535), 
        .Y(n849) );
  OAI221XL U1395 ( .A0(n544), .A1(n1103), .B0(n1097), .B1(n564), .C0(n565), 
        .Y(n862) );
  OAI21XL U1396 ( .A0(n566), .A1(n522), .B0(cs[2]), .Y(n565) );
  CLKINVX1 U1397 ( .A(n567), .Y(n1103) );
  OAI221XL U1398 ( .A0(int_i[0]), .A1(n531), .B0(n260), .B1(n532), .C0(n488), 
        .Y(n848) );
  NOR3X1 U1399 ( .A(cs[1]), .B(cs[2]), .C(cs[0]), .Y(n539) );
  XNOR2X1 U1400 ( .A(tmp_T0[3]), .B(n277), .Y(n343) );
  XNOR2X1 U1401 ( .A(tmp_T0[0]), .B(n1152), .Y(n346) );
  XNOR2X1 U1402 ( .A(tmp_T0[1]), .B(n1151), .Y(n345) );
  XNOR2X1 U1403 ( .A(tmp_T0[2]), .B(n1150), .Y(n344) );
  OAI211X1 U1404 ( .A0(n347), .A1(n268), .B0(n379), .C0(n380), .Y(n741) );
  AOI2BB2X1 U1405 ( .B0(\Tree_1[2][0] ), .B1(n352), .A0N(n353), .A1N(n264), 
        .Y(n379) );
  AOI222XL U1406 ( .A0(tmp_T1[0]), .A1(n1002), .B0(\Tree_1[4][0] ), .B1(n1008), 
        .C0(\Tree_1[1][0] ), .C1(n351), .Y(n380) );
  OAI211X1 U1407 ( .A0(n347), .A1(n276), .B0(n367), .C0(n368), .Y(n725) );
  AOI222XL U1408 ( .A0(tmp_T0[0]), .A1(n1002), .B0(\Tree_0[4][0] ), .B1(n1008), 
        .C0(\Tree_0[1][0] ), .C1(n351), .Y(n368) );
  OAI211X1 U1409 ( .A0(n347), .A1(n266), .B0(n373), .C0(n374), .Y(n733) );
  AOI222XL U1410 ( .A0(tmp_T1[2]), .A1(n1002), .B0(\Tree_1[4][2] ), .B1(n1008), 
        .C0(\Tree_1[1][2] ), .C1(n351), .Y(n374) );
  OAI211X1 U1411 ( .A0(n347), .A1(n274), .B0(n361), .C0(n362), .Y(n717) );
  AOI222XL U1412 ( .A0(tmp_T0[2]), .A1(n1002), .B0(\Tree_0[4][2] ), .B1(n1008), 
        .C0(\Tree_0[1][2] ), .C1(n351), .Y(n362) );
  OAI211X1 U1413 ( .A0(n347), .A1(n265), .B0(n370), .C0(n371), .Y(n729) );
  AOI222XL U1414 ( .A0(tmp_T1[3]), .A1(n1002), .B0(\Tree_1[4][3] ), .B1(n1008), 
        .C0(\Tree_1[1][3] ), .C1(n351), .Y(n371) );
  OAI211X1 U1415 ( .A0(n347), .A1(n273), .B0(n348), .C0(n349), .Y(n713) );
  AOI222XL U1416 ( .A0(tmp_T0[3]), .A1(n1002), .B0(\Tree_0[4][3] ), .B1(n1008), 
        .C0(\Tree_0[1][3] ), .C1(n351), .Y(n349) );
  OAI211X1 U1417 ( .A0(n347), .A1(n267), .B0(n376), .C0(n377), .Y(n737) );
  AOI222XL U1418 ( .A0(tmp_T1[1]), .A1(n1002), .B0(\Tree_1[4][1] ), .B1(n1008), 
        .C0(\Tree_1[1][1] ), .C1(n351), .Y(n377) );
  OAI211X1 U1419 ( .A0(n347), .A1(n275), .B0(n364), .C0(n365), .Y(n721) );
  AOI222XL U1420 ( .A0(tmp_T0[1]), .A1(n1002), .B0(\Tree_0[4][1] ), .B1(n1008), 
        .C0(\Tree_0[1][1] ), .C1(n351), .Y(n365) );
  OAI211X1 U1421 ( .A0(n533), .A1(n1107), .B0(n556), .C0(n557), .Y(n858) );
  CLKINVX1 U1422 ( .A(n561), .Y(n1107) );
  AOI21X1 U1423 ( .A0(int_j[2]), .A1(n558), .B0(n536), .Y(n557) );
  OAI21XL U1424 ( .A0(n1088), .A1(n251), .B0(n534), .Y(n558) );
  NAND3X1 U1425 ( .A(n255), .B(n253), .C(N488), .Y(n544) );
  AND3X2 U1426 ( .A(n1104), .B(n255), .C(n387), .Y(n1023) );
  NOR3X1 U1427 ( .A(n458), .B(cnt2[0]), .C(n150), .Y(n546) );
  OAI22XL U1428 ( .A0(n986), .A1(n295), .B0(n1050), .B1(n296), .Y(n704) );
  OAI22XL U1429 ( .A0(n986), .A1(n289), .B0(n1049), .B1(n290), .Y(n662) );
  OAI22XL U1430 ( .A0(n986), .A1(n290), .B0(n1049), .B1(n291), .Y(n669) );
  OAI22XL U1431 ( .A0(n986), .A1(n291), .B0(n1049), .B1(n292), .Y(n676) );
  OAI22XL U1432 ( .A0(n986), .A1(n292), .B0(n1049), .B1(n293), .Y(n683) );
  OAI22XL U1433 ( .A0(n986), .A1(n293), .B0(n1049), .B1(n294), .Y(n690) );
  OAI22XL U1434 ( .A0(n986), .A1(n294), .B0(n1049), .B1(n295), .Y(n697) );
  OAI2BB2XL U1435 ( .B0(n545), .B1(n150), .A0N(n545), .A1N(cnt2[0]), .Y(n853)
         );
  OAI22XL U1436 ( .A0(n529), .A1(n259), .B0(int_i[1]), .B1(n530), .Y(n847) );
  OAI22XL U1437 ( .A0(n545), .A1(n151), .B0(cnt2[0]), .B1(n1096), .Y(n852) );
  AND2XL U1438 ( .A(n577), .B(n1010), .Y(n578) );
  OAI22XL U1439 ( .A0(n1049), .A1(n298), .B0(n297), .B1(n986), .Y(n649) );
  OAI22XL U1440 ( .A0(n298), .A1(n986), .B0(n1049), .B1(n299), .Y(n650) );
  OAI22XL U1441 ( .A0(n986), .A1(n299), .B0(n1049), .B1(n300), .Y(n651) );
  OAI22XL U1442 ( .A0(n986), .A1(n300), .B0(n1049), .B1(n301), .Y(n652) );
  OAI22XL U1443 ( .A0(n986), .A1(n301), .B0(n1049), .B1(n302), .Y(n653) );
  OAI22XL U1444 ( .A0(n986), .A1(n302), .B0(n1049), .B1(n303), .Y(n654) );
  OAI22XL U1445 ( .A0(n986), .A1(n303), .B0(n1049), .B1(n304), .Y(n655) );
  OAI22XL U1446 ( .A0(n277), .A1(n328), .B0(n1111), .B1(n1050), .Y(n645) );
  OAI21XL U1447 ( .A0(n255), .A1(n559), .B0(n524), .Y(n860) );
  OAI21XL U1495 ( .A0(n986), .A1(n296), .B0(n1050), .Y(n712) );
  OAI2BB2XL U1497 ( .B0(n1051), .B1(n281), .A0N(HC1[7]), .A1N(n1052), .Y(n643)
         );
  OAI2BB2XL U1499 ( .B0(n1055), .B1(n281), .A0N(HC3[7]), .A1N(n1056), .Y(n641)
         );
  OAI2BB2XL U1500 ( .B0(n1057), .B1(n281), .A0N(HC4[7]), .A1N(n1058), .Y(n640)
         );
  OAI2BB2XL U1501 ( .B0(n1059), .B1(n281), .A0N(HC5[7]), .A1N(n1060), .Y(n639)
         );
  OAI2BB2XL U1509 ( .B0(n1051), .B1(n284), .A0N(HC1[4]), .A1N(n1052), .Y(n608)
         );
  OAI2BB2XL U1511 ( .B0(n1055), .B1(n284), .A0N(HC3[4]), .A1N(n1056), .Y(n606)
         );
  OAI2BB2XL U1512 ( .B0(n1057), .B1(n284), .A0N(HC4[4]), .A1N(n1058), .Y(n605)
         );
  OAI2BB2XL U1513 ( .B0(n1059), .B1(n284), .A0N(HC5[4]), .A1N(n1060), .Y(n604)
         );
  OAI2BB2XL U1515 ( .B0(n1051), .B1(n285), .A0N(HC1[3]), .A1N(n1052), .Y(n615)
         );
  OAI2BB2XL U1517 ( .B0(n1055), .B1(n285), .A0N(HC3[3]), .A1N(n1056), .Y(n613)
         );
  OAI2BB2XL U1518 ( .B0(n1057), .B1(n285), .A0N(HC4[3]), .A1N(n1058), .Y(n612)
         );
  OAI2BB2XL U1519 ( .B0(n1059), .B1(n285), .A0N(HC5[3]), .A1N(n1060), .Y(n611)
         );
  OAI2BB2XL U1521 ( .B0(n1051), .B1(n286), .A0N(HC1[2]), .A1N(n1052), .Y(n622)
         );
  OAI2BB2XL U1523 ( .B0(n1055), .B1(n286), .A0N(HC3[2]), .A1N(n1056), .Y(n620)
         );
  OAI2BB2XL U1524 ( .B0(n1057), .B1(n286), .A0N(HC4[2]), .A1N(n1058), .Y(n619)
         );
  OAI2BB2XL U1525 ( .B0(n1059), .B1(n286), .A0N(HC5[2]), .A1N(n1060), .Y(n618)
         );
  OAI2BB2XL U1527 ( .B0(n1051), .B1(n287), .A0N(HC1[1]), .A1N(n1052), .Y(n629)
         );
  OAI2BB2XL U1529 ( .B0(n1055), .B1(n287), .A0N(HC3[1]), .A1N(n1056), .Y(n627)
         );
  OAI2BB2XL U1530 ( .B0(n1057), .B1(n287), .A0N(HC4[1]), .A1N(n1058), .Y(n626)
         );
  OAI2BB2XL U1531 ( .B0(n1059), .B1(n287), .A0N(HC5[1]), .A1N(n1060), .Y(n625)
         );
  OAI2BB2XL U1532 ( .B0(n1061), .B1(n287), .A0N(HC6[1]), .A1N(n1062), .Y(n624)
         );
  OAI2BB2XL U1533 ( .B0(n1051), .B1(n288), .A0N(HC1[0]), .A1N(n1052), .Y(n636)
         );
  OAI2BB2XL U1535 ( .B0(n1055), .B1(n288), .A0N(HC3[0]), .A1N(n1056), .Y(n634)
         );
  OAI2BB2XL U1536 ( .B0(n1057), .B1(n288), .A0N(HC4[0]), .A1N(n1058), .Y(n633)
         );
  OAI2BB2XL U1537 ( .B0(n1059), .B1(n288), .A0N(HC5[0]), .A1N(n1060), .Y(n632)
         );
  OAI2BB2XL U1538 ( .B0(n1061), .B1(n288), .A0N(HC6[0]), .A1N(n1062), .Y(n631)
         );
  OAI2BB2XL U1539 ( .B0(n1051), .B1(n289), .A0N(M1[7]), .A1N(n1052), .Y(n661)
         );
  OAI2BB2XL U1541 ( .B0(n1055), .B1(n289), .A0N(M3[7]), .A1N(n1056), .Y(n659)
         );
  OAI2BB2XL U1542 ( .B0(n1057), .B1(n289), .A0N(M4[7]), .A1N(n1058), .Y(n658)
         );
  OAI2BB2XL U1543 ( .B0(n1059), .B1(n289), .A0N(M5[7]), .A1N(n1060), .Y(n657)
         );
  OAI2BB2XL U1544 ( .B0(n1061), .B1(n289), .A0N(M6[7]), .A1N(n1062), .Y(n656)
         );
  OAI21XL U1545 ( .A0(n253), .A1(n559), .B0(n556), .Y(n859) );
  NAND4X1 U1546 ( .A(n552), .B(n553), .C(n554), .D(n546), .Y(n551) );
  XNOR2X1 U1547 ( .A(int_j[2]), .B(int_i[2]), .Y(n554) );
  XNOR2X1 U1548 ( .A(\int_k[2] ), .B(N296), .Y(n390) );
  OAI21XL U1549 ( .A0(n986), .A1(n304), .B0(n324), .Y(n705) );
  CLKINVX1 U1550 ( .A(RegA_v[7]), .Y(n1153) );
  AND3X2 U1551 ( .A(n387), .B(N296), .C(n388), .Y(n1024) );
  CLKINVX1 U1552 ( .A(node[0]), .Y(n1152) );
  CLKINVX1 U1553 ( .A(node[1]), .Y(n1151) );
  CLKINVX1 U1554 ( .A(node[2]), .Y(n1150) );
  NOR3X2 U1555 ( .A(n310), .B(cs[0]), .C(n309), .Y(code_valid) );
  NOR2X1 U1556 ( .A(int_j[1]), .B(int_j[2]), .Y(n561) );
  NAND3X1 U1557 ( .A(n310), .B(n309), .C(cs[0]), .Y(n572) );
  OAI222XL U1558 ( .A0(n452), .A1(n984), .B0(n994), .B1(n82), .C0(n1041), .C1(
        n1162), .Y(n801) );
  OAI222XL U1559 ( .A0(n444), .A1(n984), .B0(n994), .B1(n78), .C0(n1041), .C1(
        n1193), .Y(n797) );
  OAI222XL U1560 ( .A0(n448), .A1(n984), .B0(n994), .B1(n80), .C0(n1041), .C1(
        n1178), .Y(n799) );
  OAI222XL U1561 ( .A0(n442), .A1(n984), .B0(n994), .B1(n77), .C0(n1041), .C1(
        n1200), .Y(n796) );
  OAI222XL U1562 ( .A0(n446), .A1(n984), .B0(n994), .B1(n79), .C0(n1041), .C1(
        n1186), .Y(n798) );
  OAI222XL U1563 ( .A0(n450), .A1(n984), .B0(n994), .B1(n81), .C0(n1041), .C1(
        n1170), .Y(n800) );
  OAI222XL U1564 ( .A0(n452), .A1(n991), .B0(n995), .B1(n122), .C0(n1032), 
        .C1(n1161), .Y(n793) );
  OAI222XL U1565 ( .A0(n450), .A1(n991), .B0(n995), .B1(n121), .C0(n1032), 
        .C1(n1169), .Y(n791) );
  OAI222XL U1566 ( .A0(n448), .A1(n991), .B0(n995), .B1(n120), .C0(n1032), 
        .C1(n1177), .Y(n789) );
  OAI222XL U1567 ( .A0(n446), .A1(n991), .B0(n995), .B1(n119), .C0(n1032), 
        .C1(n1185), .Y(n787) );
  OAI222XL U1568 ( .A0(n444), .A1(n991), .B0(n995), .B1(n118), .C0(n1032), 
        .C1(n1192), .Y(n785) );
  OAI222XL U1569 ( .A0(n442), .A1(n991), .B0(n995), .B1(n117), .C0(n1032), 
        .C1(n1199), .Y(n783) );
  OAI222XL U1570 ( .A0(n440), .A1(n991), .B0(n995), .B1(n116), .C0(n1032), 
        .C1(n1207), .Y(n781) );
  OAI222XL U1571 ( .A0(n453), .A1(n991), .B0(n995), .B1(n115), .C0(n1032), 
        .C1(n1159), .Y(n843) );
  OAI222XL U1572 ( .A0(n440), .A1(n997), .B0(n998), .B1(n108), .C0(n1038), 
        .C1(n1212), .Y(n827) );
  OAI222XL U1573 ( .A0(n453), .A1(n997), .B0(n998), .B1(n107), .C0(n1038), 
        .C1(n1158), .Y(n826) );
  OAI222XL U1574 ( .A0(n440), .A1(n984), .B0(n994), .B1(n76), .C0(n1041), .C1(
        n1208), .Y(n795) );
  CLKINVX12 U1575 ( .A(n1063), .Y(n1071) );
  MXI2X4 U1576 ( .A(n115), .B(n1064), .S0(n1071), .Y(n865) );
  MXI2X4 U1577 ( .A(n116), .B(n1065), .S0(n1071), .Y(n866) );
  MXI2X4 U1578 ( .A(n117), .B(n1066), .S0(n1071), .Y(n867) );
  MXI2X4 U1579 ( .A(n118), .B(n1067), .S0(n1071), .Y(n868) );
  MXI2X4 U1580 ( .A(n119), .B(n1068), .S0(n1071), .Y(n869) );
  MXI2X4 U1581 ( .A(n120), .B(n1069), .S0(n1071), .Y(n870) );
  MXI2X4 U1582 ( .A(n121), .B(n1070), .S0(n1071), .Y(n871) );
  MXI2X4 U1583 ( .A(n122), .B(n1072), .S0(n1071), .Y(n872) );
  MXI2X4 U1584 ( .A(n75), .B(n1076), .S0(n1030), .Y(n905) );
  MXI2X4 U1585 ( .A(n76), .B(n1077), .S0(n1030), .Y(n906) );
  MXI2X4 U1586 ( .A(n77), .B(n1078), .S0(n1030), .Y(n907) );
  MXI2X4 U1587 ( .A(n78), .B(n1079), .S0(n1030), .Y(n908) );
  MXI2X4 U1588 ( .A(n79), .B(n1080), .S0(n1030), .Y(n909) );
  MXI2X4 U1589 ( .A(n80), .B(n1081), .S0(n1030), .Y(n910) );
  MXI2X4 U1590 ( .A(n81), .B(n1082), .S0(n1030), .Y(n911) );
  MXI2X4 U1591 ( .A(n82), .B(n1083), .S0(n1030), .Y(n912) );
  huffman_DW01_add_0 add_609 ( .A(tmp_HC), .B(addnum), .CI(1'b0), .SUM({N719, 
        N718, N717, N716, N715, N714, N713, N712}) );
  huffman_DW01_add_1 add_461 ( .A(RegA_v), .B(RegB_v), .CI(1'b0), .SUM({N499, 
        N498, N497, N496, N495, N494, N493, N492}) );
  huffman_DW01_inc_0 add_424_S2 ( .A({cnt[6:1], n1044}), .SUM({N446, N445, 
        N444, N443, N442, N441, N440}) );
  huffman_DW01_inc_1 add_411 ( .A(CNT6), .SUM({N425, N424, N423, N422, N421, 
        N420, N419, N418}) );
  huffman_DW01_inc_2 add_410 ( .A(CNT5), .SUM({N417, N416, N415, N414, N413, 
        N412, N411, N410}) );
  huffman_DW01_inc_3 add_409 ( .A(CNT4), .SUM({N409, N408, N407, N406, N405, 
        N404, N403, N402}) );
  huffman_DW01_inc_4 add_408 ( .A(CNT3), .SUM({N401, N400, N399, N398, N397, 
        N396, N395, N394}) );
  huffman_DW01_inc_5 add_407 ( .A(CNT2), .SUM({N393, N392, N391, N390, N389, 
        N388, N387, N386}) );
  huffman_DW01_inc_6 add_406 ( .A(CNT1), .SUM({N385, N384, N383, N382, N381, 
        N380, N379, N378}) );
  BUFX16 U860 ( .A(gray_valid), .Y(net7492) );
  NOR3X4 U859 ( .A(gray_data[3]), .B(gray_data[5]), .C(gray_data[4]), .Y(n933)
         );
  AND2X6 U757 ( .A(n933), .B(net5514), .Y(net7188) );
  NOR2X6 U759 ( .A(gray_data[7]), .B(gray_data[6]), .Y(net5514) );
  CLKINVX8 U857 ( .A(gray_data[2]), .Y(net7494) );
  NOR3X4 U856 ( .A(net7469), .B(net7433), .C(gray_data[1]), .Y(net5512) );
  INVX8 U855 ( .A(net7494), .Y(net7433) );
  AOI2BB2X4 U1009 ( .B0(n572), .B1(net5697), .A0N(net5697), .A1N(n539), .Y(
        n569) );
  NAND2X6 U761 ( .A(n938), .B(net5697), .Y(n935) );
  BUFX16 U854 ( .A(gray_valid), .Y(net5697) );
  NOR3X8 U853 ( .A(net5701), .B(net5501), .C(net7385), .Y(net5500) );
  NOR3X8 U850 ( .A(gray_data[3]), .B(gray_data[5]), .C(gray_data[4]), .Y(n932)
         );
  NAND2X8 U758 ( .A(net5514), .B(n932), .Y(net7388) );
  CLKINVX12 U849 ( .A(net7388), .Y(net7189) );
  NAND2X8 U848 ( .A(net7189), .B(net5488), .Y(net7366) );
  CLKMX2X4 U846 ( .A(CNT3[7]), .B(N401), .S0(net5660), .Y(n881) );
  DFFX1 \tmp_MK_reg[0]  ( .D(n712), .CK(clk), .Q(n1243), .QN(n296) );
  DFFX1 \tmp_MK_reg[1]  ( .D(n704), .CK(clk), .Q(n1242), .QN(n295) );
  DFFX1 \tmp_MK_reg[6]  ( .D(n669), .CK(clk), .Q(n1241), .QN(n290) );
  DFFX1 \tmp_MK_reg[5]  ( .D(n676), .CK(clk), .Q(n1240), .QN(n291) );
  DFFX1 \tmp_MK_reg[4]  ( .D(n683), .CK(clk), .Q(n1239), .QN(n292) );
  DFFX1 \tmp_MK_reg[3]  ( .D(n690), .CK(clk), .Q(n1238), .QN(n293) );
  DFFX1 \tmp_MK_reg[2]  ( .D(n697), .CK(clk), .Q(n1237), .QN(n294) );
  EDFFHQX1 \HC3_reg[6]  ( .D(tmp_HC[6]), .E(n1234), .CK(clk), .Q(n1246) );
  EDFFHQX1 \HC6_reg[6]  ( .D(tmp_HC[6]), .E(n1233), .CK(clk), .Q(n1251) );
  EDFFHQX1 \HC4_reg[5]  ( .D(tmp_HC[5]), .E(n1235), .CK(clk), .Q(n1248) );
  EDFFHQX1 \HC3_reg[5]  ( .D(tmp_HC[5]), .E(n1234), .CK(clk), .Q(n1247) );
  EDFFHQX1 \HC1_reg[6]  ( .D(tmp_HC[6]), .E(n1232), .CK(clk), .Q(n1244) );
  EDFFHQX1 \HC1_reg[5]  ( .D(tmp_HC[5]), .E(n1232), .CK(clk), .Q(n1245) );
  EDFFHQX1 \HC5_reg[6]  ( .D(tmp_HC[6]), .E(n1231), .CK(clk), .Q(n1249) );
  EDFFHQX1 \HC5_reg[5]  ( .D(tmp_HC[5]), .E(n1231), .CK(clk), .Q(n1250) );
  DFFXL \RegA_t_reg[3]  ( .D(n773), .CK(clk), .Q(RegA_t[3]), .QN(n1127) );
  DFFXL \RegA_t_reg[0]  ( .D(n776), .CK(clk), .Q(RegA_t[0]), .QN(n1142) );
  DFFXL \ListB_reg[0][7]  ( .D(n843), .CK(clk), .Q(\ListB[0][7] ), .QN(n1159)
         );
  DFFXL \ListB_reg[0][6]  ( .D(n781), .CK(clk), .Q(\ListB[0][6] ), .QN(n1207)
         );
  DFFXL \ListB_reg[0][5]  ( .D(n783), .CK(clk), .Q(\ListB[0][5] ), .QN(n1199)
         );
  DFFXL \ListB_reg[0][4]  ( .D(n785), .CK(clk), .Q(\ListB[0][4] ), .QN(n1192)
         );
  DFFXL \ListB_reg[0][3]  ( .D(n787), .CK(clk), .Q(\ListB[0][3] ), .QN(n1185)
         );
  DFFXL \ListB_reg[0][2]  ( .D(n789), .CK(clk), .Q(\ListB[0][2] ), .QN(n1177)
         );
  DFFXL \ListB_reg[0][1]  ( .D(n791), .CK(clk), .Q(\ListB[0][1] ), .QN(n1169)
         );
  DFFXL \ListB_reg[0][0]  ( .D(n793), .CK(clk), .Q(\ListB[0][0] ), .QN(n1161)
         );
  EDFFHQX2 \HC2_reg[4]  ( .D(tmp_HC[4]), .E(n1236), .CK(clk), .Q(HC2[4]) );
  EDFFHQX2 \HC2_reg[3]  ( .D(tmp_HC[3]), .E(n1236), .CK(clk), .Q(HC2[3]) );
  EDFFHQX2 \HC2_reg[2]  ( .D(tmp_HC[2]), .E(n1236), .CK(clk), .Q(HC2[2]) );
  EDFFHQX2 \HC2_reg[1]  ( .D(tmp_HC[1]), .E(n1236), .CK(clk), .Q(HC2[1]) );
  EDFFHQX2 \HC2_reg[0]  ( .D(tmp_HC[0]), .E(n1236), .CK(clk), .Q(HC2[0]) );
  EDFFHQX2 \M2_reg[7]  ( .D(n1017), .E(n1236), .CK(clk), .Q(M2[7]) );
  DFFRX2 \int_k_reg[1]  ( .D(n860), .CK(clk), .RN(n1084), .Q(N296), .QN(n255)
         );
  EDFFHQX2 \HC2_reg[6]  ( .D(tmp_HC[6]), .E(n1236), .CK(clk), .Q(HC2[6]) );
  EDFFHQX2 \HC2_reg[5]  ( .D(tmp_HC[5]), .E(n1236), .CK(clk), .Q(HC2[5]) );
  EDFFHQX2 \HC4_reg[6]  ( .D(tmp_HC[6]), .E(n1235), .CK(clk), .Q(HC4[6]) );
  EDFFHQX2 \HC6_reg[5]  ( .D(tmp_HC[5]), .E(n1233), .CK(clk), .Q(HC6[5]) );
  EDFFHQX2 \M2_reg[0]  ( .D(n1243), .E(n1236), .CK(clk), .Q(M2[0]) );
  EDFFHQX2 \M6_reg[0]  ( .D(n1243), .E(n1233), .CK(clk), .Q(M6[0]) );
  EDFFHQX2 \M4_reg[0]  ( .D(n1243), .E(n1235), .CK(clk), .Q(M4[0]) );
  EDFFHQX2 \M3_reg[0]  ( .D(n1243), .E(n1234), .CK(clk), .Q(M3[0]) );
  EDFFHQX2 \M1_reg[0]  ( .D(n1243), .E(n1232), .CK(clk), .Q(M1[0]) );
  EDFFHQX2 \M5_reg[0]  ( .D(n1243), .E(n1231), .CK(clk), .Q(M5[0]) );
  EDFFHQX2 \M2_reg[6]  ( .D(n1241), .E(n1236), .CK(clk), .Q(M2[6]) );
  EDFFHQX2 \M2_reg[5]  ( .D(n1240), .E(n1236), .CK(clk), .Q(M2[5]) );
  EDFFHQX2 \M2_reg[4]  ( .D(n1239), .E(n1236), .CK(clk), .Q(M2[4]) );
  EDFFHQX2 \M2_reg[3]  ( .D(n1238), .E(n1236), .CK(clk), .Q(M2[3]) );
  EDFFHQX2 \M2_reg[2]  ( .D(n1237), .E(n1236), .CK(clk), .Q(M2[2]) );
  EDFFHQX2 \M2_reg[1]  ( .D(n1242), .E(n1236), .CK(clk), .Q(M2[1]) );
  EDFFHQX2 \M6_reg[6]  ( .D(n1241), .E(n1233), .CK(clk), .Q(M6[6]) );
  EDFFHQX2 \M6_reg[5]  ( .D(n1240), .E(n1233), .CK(clk), .Q(M6[5]) );
  EDFFHQX2 \M6_reg[4]  ( .D(n1239), .E(n1233), .CK(clk), .Q(M6[4]) );
  EDFFHQX2 \M4_reg[6]  ( .D(n1241), .E(n1235), .CK(clk), .Q(M4[6]) );
  EDFFHQX2 \M4_reg[5]  ( .D(n1240), .E(n1235), .CK(clk), .Q(M4[5]) );
  EDFFHQX2 \M4_reg[4]  ( .D(n1239), .E(n1235), .CK(clk), .Q(M4[4]) );
  EDFFHQX2 \M4_reg[3]  ( .D(n1238), .E(n1235), .CK(clk), .Q(M4[3]) );
  EDFFHQX2 \M3_reg[6]  ( .D(n1241), .E(n1234), .CK(clk), .Q(M3[6]) );
  EDFFHQX2 \M3_reg[5]  ( .D(n1240), .E(n1234), .CK(clk), .Q(M3[5]) );
  EDFFHQX2 \M3_reg[4]  ( .D(n1239), .E(n1234), .CK(clk), .Q(M3[4]) );
  EDFFHQX2 \M3_reg[3]  ( .D(n1238), .E(n1234), .CK(clk), .Q(M3[3]) );
  EDFFHQX2 \M6_reg[3]  ( .D(n1238), .E(n1233), .CK(clk), .Q(M6[3]) );
  EDFFHQX2 \M6_reg[2]  ( .D(n1237), .E(n1233), .CK(clk), .Q(M6[2]) );
  EDFFHQX2 \M6_reg[1]  ( .D(n1242), .E(n1233), .CK(clk), .Q(M6[1]) );
  EDFFHQX2 \M4_reg[2]  ( .D(n1237), .E(n1235), .CK(clk), .Q(M4[2]) );
  EDFFHQX2 \M4_reg[1]  ( .D(n1242), .E(n1235), .CK(clk), .Q(M4[1]) );
  EDFFHQX2 \M3_reg[2]  ( .D(n1237), .E(n1234), .CK(clk), .Q(M3[2]) );
  EDFFHQX2 \M3_reg[1]  ( .D(n1242), .E(n1234), .CK(clk), .Q(M3[1]) );
  EDFFHQX2 \M1_reg[6]  ( .D(n1241), .E(n1232), .CK(clk), .Q(M1[6]) );
  EDFFHQX2 \M1_reg[5]  ( .D(n1240), .E(n1232), .CK(clk), .Q(M1[5]) );
  EDFFHQX2 \M1_reg[4]  ( .D(n1239), .E(n1232), .CK(clk), .Q(M1[4]) );
  EDFFHQX2 \M1_reg[3]  ( .D(n1238), .E(n1232), .CK(clk), .Q(M1[3]) );
  EDFFHQX2 \M1_reg[2]  ( .D(n1237), .E(n1232), .CK(clk), .Q(M1[2]) );
  EDFFHQX2 \M1_reg[1]  ( .D(n1242), .E(n1232), .CK(clk), .Q(M1[1]) );
  EDFFHQX2 \M5_reg[6]  ( .D(n1241), .E(n1231), .CK(clk), .Q(M5[6]) );
  EDFFHQX2 \M5_reg[5]  ( .D(n1240), .E(n1231), .CK(clk), .Q(M5[5]) );
  EDFFHQX2 \M5_reg[4]  ( .D(n1239), .E(n1231), .CK(clk), .Q(M5[4]) );
  EDFFHQX2 \M5_reg[3]  ( .D(n1238), .E(n1231), .CK(clk), .Q(M5[3]) );
  EDFFHQX2 \HC2_reg[7]  ( .D(tmp_HC[7]), .E(n1236), .CK(clk), .Q(HC2[7]) );
  EDFFHQX2 \M5_reg[2]  ( .D(n1237), .E(n1231), .CK(clk), .Q(M5[2]) );
  EDFFHQX2 \M5_reg[1]  ( .D(n1242), .E(n1231), .CK(clk), .Q(M5[1]) );
  EDFFHQX2 \HC6_reg[7]  ( .D(tmp_HC[7]), .E(n1233), .CK(clk), .Q(HC6[7]) );
  EDFFHQX2 \HC6_reg[4]  ( .D(tmp_HC[4]), .E(n1233), .CK(clk), .Q(HC6[4]) );
  EDFFHQX2 \HC6_reg[3]  ( .D(tmp_HC[3]), .E(n1233), .CK(clk), .Q(HC6[3]) );
  EDFFHQX2 \HC6_reg[2]  ( .D(tmp_HC[2]), .E(n1233), .CK(clk), .Q(HC6[2]) );
  NOR3X8 U747 ( .A(n931), .B(net7433), .C(net7385), .Y(net5488) );
  NAND2X4 U807 ( .A(gray_data[0]), .B(gray_data[1]), .Y(n931) );
  CLKINVX16 U812 ( .A(n940), .Y(n1009) );
  CLKINVX16 U847 ( .A(net7366), .Y(net5660) );
  NAND2X8 U851 ( .A(net7189), .B(net5512), .Y(n1063) );
  CLKBUFX6 U852 ( .A(n393), .Y(n1032) );
  CLKMX2X4 U858 ( .A(CNT5[3]), .B(N413), .S0(net5661), .Y(n893) );
  CLKMX2X4 U861 ( .A(CNT5[2]), .B(N412), .S0(net5661), .Y(n894) );
  NAND2X4 U865 ( .A(gray_data[0]), .B(gray_data[2]), .Y(net5477) );
  BUFX8 U867 ( .A(gray_data[0]), .Y(net5701) );
  NAND2X6 U868 ( .A(net5475), .B(net7188), .Y(n941) );
  NOR3X6 U876 ( .A(net7390), .B(net5477), .C(net7476), .Y(net5475) );
  CLKMX2X4 U889 ( .A(CNT5[1]), .B(N411), .S0(net5661), .Y(n895) );
  INVXL U898 ( .A(n1250), .Y(n1215) );
  INVX3 U899 ( .A(n1215), .Y(HC5[5]) );
  INVXL U900 ( .A(n1249), .Y(n1217) );
  INVX3 U961 ( .A(n1217), .Y(HC5[6]) );
  INVXL U1071 ( .A(n1245), .Y(n1219) );
  INVX3 U1094 ( .A(n1219), .Y(HC1[5]) );
  INVXL U1167 ( .A(n1244), .Y(n1221) );
  INVX3 U1169 ( .A(n1221), .Y(HC1[6]) );
  INVXL U1171 ( .A(n1247), .Y(n1223) );
  INVX3 U1173 ( .A(n1223), .Y(HC3[5]) );
  INVXL U1175 ( .A(n1248), .Y(n1225) );
  INVX3 U1177 ( .A(n1225), .Y(HC4[5]) );
  INVXL U1178 ( .A(n1251), .Y(n1227) );
  INVX3 U1179 ( .A(n1227), .Y(HC6[6]) );
  INVX3 U1448 ( .A(n1061), .Y(n1233) );
  INVXL U1449 ( .A(n1246), .Y(n1229) );
  INVX3 U1450 ( .A(n1229), .Y(HC3[6]) );
  INVX3 U1451 ( .A(n315), .Y(n1235) );
  INVX3 U1452 ( .A(n318), .Y(n1232) );
  INVX3 U1453 ( .A(n314), .Y(n1231) );
  INVX3 U1454 ( .A(n316), .Y(n1234) );
  INVX3 U1455 ( .A(n317), .Y(n1236) );
  NAND2X8 U1456 ( .A(net7189), .B(n936), .Y(n934) );
  INVX12 U1457 ( .A(net5697), .Y(net7385) );
endmodule

